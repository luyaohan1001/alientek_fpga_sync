module cmos_driver(
    input           clk  ,          //配置驱动时钟
    input           rst_n,          //复位信号
    input           cmos_start,     //SDRAM初始化完成
    //摄像头接口                          
    input           cam_pclk  ,          
    input           cam_vsync ,         
    input           cam_href  ,        
    input  [7:0]    cam_data  ,       
    input  [9:0]    pixel_xpos,
    
        
    output          cmos_frame_vsync ,  
    output          cmos_frame_href  , 
    output          cmos_frame_valid , 
    output [15:0]   cmos_frame_data  ,
    output          cam_scl          , 
    output          cam_sda          ,
    output          cam_rst_n        ,  //cmos 复位信号，低电平有效
    output          cam_pwdn            //cmos 电源休眠模式选择信号
    ); 

//parameter define
parameter  SLAVE_ADDR = 7'h3c         ;  //OV5640的器件地址7'h3c
parameter  BIT_CTRL   = 1'b1          ;  //OV5640的字节地址为16位  0:8位 1:16位
parameter  CLK_FREQ   = 26'd65_000_000;  //i2c_dri模块的驱动时钟频率 65MHz
parameter  I2C_FREQ   = 18'd250_000   ;  //I2C的SCL时钟频率,不超过400KHz
parameter  CMOS_H_PIXEL = 24'd512     ;  //CMOS水平方向像素个数,用于设置SDRAM缓存大小
parameter  CMOS_V_PIXEL = 24'd768     ;  //CMOS垂直方向像素个数,用于设置SDRAM缓存大小
    
//wire define 
wire          i2c_dri_clk;  //IIC驱动时钟
wire          i2c_done   ;  //IIC写完成
wire          i2c_exec   ;  //IIC配置完成
wire          clk_65m;      //65mhz时钟,提供给IIC驱动时钟和vga驱动时钟
wire [23:0]   i2c_data  ;   //I2C要配置的地址与数据(高8位地址,低8位数据)
wire          cam_init_done;//摄像头初始化完成
wire          sys_init_done;//系统初始化完成标志
//系统初始化完成：SDRAM和摄像头都初始化完成
//避免了在SDRAM初始化过程中向里面写入数据 
assign sys_init_done = cmos_start & cam_init_done;
//不对摄像头硬件复位,固定高电平
assign  cam_rst_n = 1'b1;
//电源休眠模式选择 0：正常模式 1：电源休眠模式
assign  cam_pwdn = 1'b0;

//I2C配置模块
i2c_ov5640_rgb565_cfg 
   #(
     .CMOS_H_PIXEL      (CMOS_H_PIXEL),
     .CMOS_V_PIXEL      (CMOS_V_PIXEL)
    )   
   u_i2c_cfg(   
    .clk                (i2c_dri_clk),
    .rst_n              (rst_n),
    .i2c_done           (i2c_done),
    .i2c_exec           (i2c_exec),
    .i2c_data           (i2c_data),
    .init_done          (cam_init_done)
    );    

//I2C驱动模块
i2c_dri 
   #(
    .SLAVE_ADDR         (SLAVE_ADDR),       //参数传递
    .CLK_FREQ           (CLK_FREQ  ),              
    .I2C_FREQ           (I2C_FREQ  )                
    )   
   u_i2c_dri(   
    .clk                (clk   ),
    .rst_n              (rst_n     ),   
        
    .i2c_exec           (i2c_exec  ),   
    .bit_ctrl           (BIT_CTRL  ),   
    .i2c_rh_wl          (1'b0),             //固定为0，只用到了IIC驱动的写操作   
    .i2c_addr           (i2c_data[23:8]),   
    .i2c_data_w         (i2c_data[7:0]),   
    .i2c_data_r         (),   
    .i2c_done           (i2c_done  ),   
    .scl                (cam_scl   ),   
    .sda                (cam_sda   ),   
        
    .dri_clk            (i2c_dri_clk)       //I2C操作时钟
);    
    
//CMOS图像数据采集模块
cmos_capture_data u_cmos_capture_data(      //系统初始化完成之后再开始采集数据 
    .rst_n              (rst_n & sys_init_done), 
        
    .cam_pclk           (cam_pclk),
    .cam_vsync          (cam_vsync),
    .cam_href           (cam_href),
    .cam_data           (cam_data),
        
        
    .cmos_frame_vsync   (),
    .cmos_frame_href    (),
    .cmos_frame_valid   (cmos_frame_valid),       //数据有效使能信号
    .cmos_frame_data    (cmos_frame_data)         //有效数据 
    );
    
endmodule
