��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ����{��=B��6WD�Z.�/3����V����� ;�"5F�� 2���BKG�Y�`�'�':L;{�1����t���H&�6�W5\}�k�:�r��p̫����t�)�|��m���?���IyN� �M����J�Va�D��G�k�Yn�oN�ͅ��^�h�{P�=dnb��9�l�D��g2{�]K��LnO�v-�;�-�\䘛���Ν��%��n��l�%͗1����y�g�L��e�y�����<J�����Y�T��F�HD�C)�O�h�Pç�=�I�U���$�,��SBY��,�Q�R�xi'[wި�lfUKs`��p+��2��J]Q8J�VX���[r��c�t�Y%�K�\c$�c�8~�*)f]���6uF[������?/iw(��!~����1�*oF�v"ؤU"8l�VTU_��761v%^D�_HfkbB)DvZAA�T���q�
Ӊ�!>k6���D܄#��Ϗ6ҽ4�6�7�����n+��(𥏾[��Y:���4o��G�FE���o7������M0�[V\���eT��\�d�R��*���^t��z�:�� �"xGD2����s��H��@s�+3�G-/��y@*��ɜ�Ӆr���c�"�IƇ��[�$�ewū��B��CVT}7q���e�a�P��A���f%�@�颍�����J�M�C�w9� ���C�����"�e�ԄQ(�$��7�TK Q��od92"ι�g3{_�R�Hne������<�����f���<1@�^����re�V�q>�W�A6A�YT�x��W{�^�|����j`[��]#�Mf�4��yS4YFݒ䃻��[����þ��qS)
׮��U�Mp�9��a���S<�d�i�SeދL=je���\�D�>�ۋ���D�E����񅳠���']�S~_Sy��#*��їH��I�d�t��ֶn���d;a�s)]�<<�F�����
�\�a�`����!�݉8�{�ʲ�أ��ݪ"׼ǺW�J�ƭ! �L&�|GǉG!]�øhW�^{�}���&�	9� *��O�˝�R$��P�G�%�H�Sr�=���n��^�kѪ*x& =H�)��D�� }�+B�(�W�R�oԾ6"$�1���qi֭��	vD���J��ڳ��n�*������N8kh�}B��?
��U��d�D�&Ø�}3���A�eO��0�T)2X�5	�������}��-w!H��5\*��.��*�z�PNN���74��@��-��K��Ě�>�<
�c�&���>�*���!H�(jn���'EVBV43Ѯ��v���L��ͭ5��!�R��j�FaC_G*m��w@��TL�~T���~��%dQ���γ��R+dt2��I R��%�c)����ĉ"�,H�x%d�z{�#!{�2ȳ�·E>/�/X�(dt[�3�()����Q��h�P@<��|EI�e�ff�9檣�˅�\�xr2w�:���n1H�Կ�S; V2�'�4J��ظ�e<�,��!I�+�P���,pռ�&��%�u�d�vG-#��PWp���4�Y�B��la�g�y����ן~O��cu�zV�|]q_f~�c]�[��}L<醞�6���%v��j�=��:��(�<b�^�{�Fax��,�f��lB�� �D8����5�s�P�lhG�����2R����"BXMf�ސ4J���@0�{��tY�C�vo��FZc��H5�ze$��^��5�Qj6e�o��<�%��'&#jpAgBw���S�z\){�}����+d3C0Ԣ�r֜���p�Mj��)�O+��4�o�=�Mq	cMPމ#���	s��"(�}�^��.aw�N��k���<pf��=�}SQl	`��/w%UB:6�{��$�b��җ��]�=��� f�[��t�I$�	Rt�ci^�]��r!h�bFhQ3���t���nU7$��+�#ﴜ����/H�5��&yɳ"�G� �,��I��md#Z΢���/F���������x"�v��iBٛGK�vH����SF,�ZYl�M�K?�!�B�U�ؾ�w��ۋ�H�d �b��U�|�� Tн�Ӕ�(�U�Gٖ��)5rR�aը��i��9z�FO�T
4T'é][D�QU?��R�D�DJ��.��OF�ؘŋ�W͂<:tܫ�"R�ɵd�~>GS��u6� ���O��lL����绻�h��$C�t@z�PS�Ґ�a�$�\�lڱ5`�n���H�O�҄���R����J�>�O�� ���|>�h�����jJ��`�����0
��nl����f-s0�ӀZ �=XME}PD�ӥD�x��e�U����*��`3�J1�m���eH|Y���x�D�s$�x���z���NIO�l X���k4����\��Ic̑r��:���'�遒��|�7��Ή��y�����v���b���x���X㲷Ł�흯�~��YS����뎅ݻj@:,]]P�xS�$C��y�,�v�
+	����g��~փ��??�R|C�gF+x�BD��J/���fJ�1՚�.�#at��Av��N�;�H&���U29h��欙��b �������o�#�'D��0l𺄔��H�(�����G7i����.DH�D���91�S�z)���'f��oya6�fuR7�M����(�[�T�pG.o��wR�e�uV���Z��n��ay�+(%�@�8	�!�N"o�gXz/]딞�RA߼f_�<�D8�%N���]�R*�br_�
+KK��J"�k5pX������7�ފ��xh�|M�t�g����%�;�|�Ը��o�|�V�E��~:PR9|�\�*���T���b6�P�31�Q�h�}���c�R�e�"��Q^�{�nUKh12�"LB�p�!�F5{+����
r�Ur���c�i���MEt�u*��Ɛj($5o|�W+��/���r�)`y�O����d��>ɵocF��ا�����2JJб�j��Q��� �/)���7 �g����T	�[��R�2,��@$6�
6�XzP2i�ލ�%�8���衚=Q�d�Ͱƽ*#���^�u����K�@�op��l�e����@���<�Z�t�d!W|_<x�}�,�������3�J��eme���,���@>e\j�-������i
#M�/h�}+���ڐ�D�GR�.%�A��]�s��1��{�@F�c�<��\�bc�k�j����X�(|�+����� /k���:g��	,�c�s�%wwU�:P�����3�P�Dg�)G�K�mű��z�=:=F������B��I�5<�u�cl���C9�Q�Q2��w��[�ʁ���4��u�U	 �R;�נC߱�Ksi�u���D�XOh�[�D\�"����v[~��^ }���b�[0�{��n�f�|�x��M��]�Gҫ���"�Y��H�eG�Yy_G��΂�"��:E�bw0�g\��9���_��`�¨��s�zlHFS�"�iܡ�'osE��Ijv�Q�J�+oau�D˿Qވ��>Hs��N����@�}��q�7�X�/����xMl���)BP3��,�6
bw���?2[�0$8�����r�	a<&]%y��ŷ��T�x��ϰ����y��;��>��~���e���r���5�w\y���O�bQ�]��m/ѽ;�!�'��4����O#��w���VO��<��v�XX�kr���KHMj�E��J%`^�?p����e
�P����YX��sA-]
�q��.��tN��i���W�i��B�B�NئI̋��y�G�y^�Q��@%�}9g O�*����(8�Eob���Z�w���=�7ˤ) �B���g�h�br���e_`؄'S�1~i��q�5F��=]�Jځ�O��b�,�}S�k'I+���H��A��AQ��c?��PI���Vl�:Ĥ���	�70'A��vs%��{���*Ѳ~�@�����V˿�0s���tE�P�|����-����+JG�o7S#�D��
]=�H)&).p� ��</�����x��u��@��*Ի�����Z���MA���/�h���w�rv�@ŭ�dN��ݥ�����VU2��M[w�[<O���^���Rb��r��q�zx��m�������{g����_�?+C|�@E�T$�~�o#~b�]$�ύ������>��?��1?ڻ��z�E��p�jY����ƈG��(EC��O�UϞj��Y8�BV&�1YmƁ"#�� v_N�A���)NЇ6�����ݭᡘ�k녾}�k�u{�Ę��������6��N��K���j��y:��f9�j3�#m��V֌Hk��
�oh��ԧI|J�m�`X2_H�\.�t3�Z�R�y<X��u��p�t��<f}�	�R^8���yH��L���]LFFD�!}l�C���=�k��x�y�,M�D ��nc��)�����'�C�*��pl�U�ZZc�We;C�Ѵ��I���\�ա��Z��o'�U�몿K���h\�����d�h�(v�����0'6��-�Ǖt�0W�uV���[t素��7N���'�'ȭ
|��esS|�@~o($}"?�:Ud�|���L;�INy��LZfG��Ս��X�F�U_/O��o�_ ��u�Δ�q�N�e��g\����l��u�|hu@���H��T9U��׶��� �WRK�Cw���/b�w�D�+�^S>Зe�Ce�$�L[o�V�j�ilE���9I+�(qL�c��1DD��Hv��㟳��LK��1r8�A�߀%�M�;|�d)��թP����Z���5X�(fX1浗R�v��s��_���4yΑ��$s׷e�u@����w�V����a=C���o�_~ �������=nF���M��nI:�_0*���{
���Ƹ�FS���>Y��F*'s�����ހ=�c��;j2m\:by��K�Q�C8l�u(�f�xZ\d����Ҭ����`ƙ,���gOH�N*���V�� �O/��ro&֩f_��/w�'�i��,)� O(�	=w��~*�ֱc_�k��p]�Kj�����Tr=�7�&����|D��f�m?t�%�"��i�C9$�.�EH\�T�a:0��,ї:m�V�ǧ��5v�$p��`=%�V2���3|��YP/i<e��)��m����ug�wR1W����y�mw�}�	�g�| ��s^^�)8�8xP�ɇ� `6�?*0D���5]F�ҝn�n:`
���3N�N�ߡ��'���F0���XDO'q���%@���W���q ae�{����R���P{��Y���H�n��@�K���p씌��[��ߏ;W_�֩���4P`���R�#o��_����ΐ�Y���ڴ��LI���
�E2R�n,��iI���Ҷ٣_� u��!�F���Y7�wռ�Xj6���z���*���q���Y��qT��1��,�W�������D�u �Z�z9)��_H+��4Fv�'ǖ�I�b.r�8�-�
����Q=�[�"��"_Az�F�V�32j�/�I}�UT�jy+I����S��7Q�*�n/=xF�A"�?X�����m� ��T�9��!>���@�߰Q^͎�/�.����A�lش�\�*���z$�(��Dm����n��jI�ݭ��x�:�ף_ĶQç 6�����	���p-�7�G�]�)T
Ȁ'QX�i�Xf",�KM<�H��_�:�?\�V�6tቇ���{�\މ,
��ۯ�����T �SV2H��9�t;�qz�g%Ɖ�&��o��j)�G�,I�5�6�������V��&q���=<Q"��,��^w��75�왂p4e�4�0BNAVu�CS7�Gd!��c,�7M@��u�p�����VP9 � !���[�̼�O�h� V��2�5"���� �K��I)��Vղ�����;SE�Ӏ6��3��չ�X[#�d/�<KӸ��>�}����#�%w���������׭���T>II�,��`�4�2�b:�@�t~u䪣U@+�r����7AI����7��ӊ�[��=���]���Q��lяgҚ^�V2 !�z� �_C��+AJ���"��i���=ɼ2�9}��^q��@���sQ�!{Jghڗ�=C���<�7��BԦ��Z�c4�9 �:=�6d����訲���Ň�аɳ� 5��U�Qa�?zf����[t´ؙ�%��P�\:���ry��r�"������R�^_4j�﹁��Z�*��T�6���6�N�ۢ��H�.J^�oK������_?�;ke0*��b�J��*�\�r�6��v���.��<C�I.�����E'��4�p'��[8nQ�2D�s�m��d�؅�P��!�y���{�[ԫ�Nҵ$��?��+�{d0(�)��Lvh�H����urf��0;�sK�.���9⻱��Z:�PǺ����u���cT�!hW���]R`*4�u9�hS���^ƅi��;��8�@x�T+�^�̄V'nAe�Am�4���.	�[�E�	��X��مޟ�*	5x����&���Eť����y�UvI �B]���Oaq�#/�'b�f��G�p�$Z����>yn`ڻ���g ���L@R;t��q�� �ߑ��q7i�I��{d�G�7]k�x�fע�����7r�Pv%�̽��%���ا@�>��GA��!\2��!bzS>xL���5��4P;�˞p9�#�p4ч�� �@^n2�z�%���2}�3�6�q���3�Ss�G����S*��Z�V��x	Ky��չ�숻ͦ���ť=�"����:&��N�(1m���O��b�[p��}�y�v�r��)3�M0I"�i1| >��ԭ����W9�	1��f� X��v�䉗)2ċJ��a@�F3�tx���ɲ���a�hk�2������i�d����������ٜ76}Cؒ��>�d��h�I��e�,�[���!
 �G@ڗ����1R�÷����k�5y�c���7f����S+�T[b��R�5��q�&��R���]�[�>a)�~�d5e��=Kή��K��i`�m���'H�8�����a�w� ��WNt�&NU�)���Pu-���v�SJ-�ƅ}�F�+�Y���9;W�{��v��?v/���H�����7 ��ߛ�,�q�V��<�,�m�H�H���DM��K��Dt).p��fq�,u*��0��x�c�)uG��WDqW�L�Gtc��Z�����j��a$���U)Ѱ	���`H�5E9��������l��d��i9�g!1�x��T�6E��X��~`_Ș���"���Y�d�k����K\6�<o��;�'�����N
49��?L�����K�!�j�p#cӪ��6zDN�R���\�N�#F��"E�1E�:��m��K�n��"��oVT9�}�۶���"n�B}�v�.�ڢ��|ʺ�H�a
�.�Ũ~! ��8x '.���ū�7��,�6ce5Z��o-.��1�"�ïhC\�ҽ�~(��.�饉^]�3�cw	A��p6��ɿrݹ�0Q&��[���Wh1�ԥ��v� �6yRi������;���֐�Cix`@�l�|kU����È�%$��~�ue�����۬���g9������ZE�J�~��۸��{&ч\��ǣںS e�5���UȜ�h��l|��`�*N[��p��P�����m9�;}B� �r�w�@��a^U�YJ�i\��N[2}����(3��4:���i*6u�n�ބ�"���1�:v�k��0$�XB^6��"rc�4�x�0�hP^�Q<�+g�چ�Qrѫ q�0�s��Ƀ���>���(�f��ḶubF�_�/��#Z�>4���D�-���:ح�Ǳ;��,e�Q�&v!5� �l7�+�"ع��8	����WL���E�����^o712޷��k�*����f� ��F�����t�U�#��4bV`bM�=<�'?�{����+��j��`�9�c�����Z^?�=�(<��`�>�M&�h�WNvG>
џP{�J!؟X�8e`m@�U{� �����6Z�̾0P�K�<���s�'�=�6��E���/K{}90��j�'�u+�r�j��vy��i�ǜYAw�p�>����T�;�?g=kݤ�h*1�]W�����fy<��3d�?��<�3��ӯ��K�k���1�mg��-y_�v9s9x%��AZ���/=��U��S_���D�� ��э˓-u_��L�.�w/R�j�J����� ��61�"u�|0��8�I`|�3��P¿�/�3�jh��1����
�Wzk9��S+�NJ3��g��G[�8��:s��ԅ����A4Y�c�qk���ז�����)��H����^�� ���\���ϱ���o��ņ��.<9��yñ��P����!�o�?�!�#�΅죈���Imfh�>�G�R!���Ǒ�҇� ��@�����P�ʧ��o�7����3�߄�yHG-�D|���D�1+���|����`h��bλѹ1<��n����D�/�oKU�2���"���s�a'�zZOx�P�`��d�,TUB�9�DX7�-:���w�����N!������G�� 6/� ���V��ԴhG����YD&(K�(T��J���"��x���
E*�a�LXQ;�qt��κP!?kѾ�g=�f��y'�v!ui:@�Ej���;��2?�-��,���։�M�k�����ݍ�ERթ��ۊ��[oqj����014F>��h[�J pNr\'äL�X�jLo�	_�a�
������t��#��5��MTdBr�f|5QP���_w	��6*e�=}5���I"��mbZĜP�/�FN���m�c�I�0vGC���B0��-N��V�r�1Lb�e��^� W���;@�*�H(�a�j�]�m:�|�����T)��	7�5k[�c���)���5%�ٵK�k���]��V���^S�E�:��`C�5����E�xI7��F��s&Qi��Ɵ��y0HB;\Q�}oZ�+rTpṎ���v�;ܴ�"T�?��o罠VJ�N��^�usX�+�V� ���C5Ӧ��B�qJur����[�Sض�>�!Y5�r��$\�tP2�>3�-����A�nYJ��.��u����)�v��#֤����4ii)��cU�H����rJn ;z_[���Ү�%(��w��Y�w����g�^����P�'|����w�<��r�>z>�4��X%�G(b�=��]�mL̦a�H���: ����s�R0O+^�Ǹ�X%F��"B��~��2�)3 �Z,�Q��y�a2��~.t�Y�әr֮�a��G��hcI�Y�Z�{M���p�j=c;�<O��K8��+p����%4H��9�<ޮ\��X�]���NBޗ�%B�
��Υy8�<� �ĳMЄ�Wg|��$x�QH(E"��4� �Eb^������G���O��_ȴ�
gs���z�l�H �o|���E���B2K1`�Ql)��HYn��~��a���[��=����~σޜ}�h���n���Zbd݆t��d(�!�r�P|�%����^��b�cI����~�1X�������R� �eTD5V�|� �J�"9ݖ\� ң�
D�M��0xѼ�2���D�ɝ��x<'ˣlK���JR�2PAg��dM��Sk�����T���u�e_��=~�}1����.���"�0�K�{C�n����󕌞�&Wq�k�E[��w�[O�t�r�SM� ~�t�U?�&k�Ms����L"�}�Y/�'���ida�E.�mc(��/�S�Q=�Uo~<���k�%�׃G��- �x���n�Y �^�.�&���d��tyF��ў�pQ��5���O���Vv�(��բvO^|o�]����В�?�c���i4�E~�҂�����H��d�ǚ�*���.>������ ����Y�]�3���gov�Д��X*@������uI͸�����2[[�$|���Bl�) d�R�<���K3�u�s>F�%�
��2=��V^)���'>D����ZY��sP�bX���iړ���h lŢ�~�n{6�F�C�k��7�{4L53���g�i��ᛖ�"�iRŲ�!��1^S|��L_K��Gv3��i9���l�͈����GKf^m�yr�z5p|]�c�� ����cL�q�ƷM4�������_㪜*J�}Ni%?ԃˍM�G7�f/��=a�+?{���c�as�����!P�o_U?j��m-Nu�PТ��n��.�7uyY ��"b��1��+bx׵������a���|����+�$������(ښe)@��eȰ]-{�r�H���-4T�zr	YzH�;���;���`&�'3�*˼�3�B�G<1�! D`�Xz	��/�N��M-�f��X��D@���[$�� ��U�k=I
��=�y�|8��ߊ! ���
9V���1�s���ÍGl-a��5�L����x{�� ��ߑ����r�k�8�
*��@�4�+#fa�%=�-��/`De��:�Z���A�uxz�f`_GAZ�\GA"F������EZ� m��U���F�^ζ�^��.��h�+X�3{>�g�=���`I�7BE�
��3}���_'O�T�3��k=�����0��_���ǫ�s��5}P?�����Ȥ�"���Id�z�$�t'íN_4o,��.�,�R��JP^ ����|��2�m���#�РBv�E���r!|	�&�	�ŪI}l���	�|�
�I�5��9��C w�ο�sտ��x���Qy��Q��ќ�DGcBӫ������X�/#�ʧ���b%�w�o���~fBD�݉cֹ��`�\u�¿Uk��1C[n�A&�U�~�S�Z�5�wL���h+c-����}LB��c�O }���aN����n�pqT��H������PsH!�����`<km�=�-����&�y13
��Y��`"ƊP�]Ɯiv8��>���ۿ�_T��I����"��JFJh�Q��$S�N?���b-.!5�'�ŞD�'}��`�$+�JԳ�����P�,?�LЇ�PY��k�tp�����D��
�D	���\�b�o}�ur��l�I� ���֨(�4:��l�B�T_O���Ϸ�a�����Ƿ��C�^_�mǠ�R��dU��q_R�]�B�1B%Y����"Ǒr���BA�żbq�����n�b^'��+#�	���b�ܸ٣�1қ�{T[_��\��� ��y�juz����e$~��{�P!�G�ۘgS�s� Y�G��E�������gWK��Mq�Lxr�f�A'P@W�`57Fg5e��+��ɥ� ���^ʑL:� ݞѻ��>g���.T)��o��?�"Sw�&8f;��u)2���O^+��ӈ��r���yi�n������c�8���K�h+���;��쭀�dD����R���J���� ��䋏��+��7��� ȱ��/@HΛ�4o�ձ���W�F��4@��"_<��S�q�d�Q@;Df	5�j}"�[ID�M���
�q���I�ztC)�}rU�^x,��V�Z]��~VӖ�S1D`�Վ�(H5a�Bd&2l�p��vl�o;�;'�8���2s����W��`�)����Ä4�W
Q4ɠ\}CXŹ1TZ�xr�u�t"j�4�֚L>�;���]��֣,H ��Mx_�r�/w����5�;"�����O�+��6��9ʋ���Z*KzqŶ�~�,kBut�!=]S.�|&��QHlt��/E���`�[i;ǉ��G��
�Q����1��{�7<��u5=j\v}Q�k��J��b�
���h�W"��aӀ����)O�b���.�����r��v81`�~yq��h��hT>m1��ƵmC�D��p�|:��2�+`�GR�"�g��Gsc?�L�BST�$!�sV�rA���й���s\���e�k�j
z���T3�d�(��y8Maj�B>r��I�������ku�d��=gw�QU��ce�{e(��_�R�q���UT[z�P%d��a�����J�P7K��JL�mj��W�=�MQ�ƄԷ`^ם�V. _��T+y��Mw��	��N�K	&�q*�r��U7���Ä&q���r�x��B����E�I�NS��abNc�����l�j+�W��](�u26ig�Y��H�ƅ�k�*�i�\���^���/8n̠AR!���Cp��$�C�ɰ6��WХ �Jc��-�q�����ͪt�����j���}츊�a�� �oI!���R��9[R<#+�{�j��$���x��Ey��
�#����5G�C]�r�����Vj0�d��(=��?מ��}@�E���˝oL3�fK���k�C��rcƵ�Nt�z��sB?ǆ�'c9�
��ۯ>p4 `|t1�OQK�i���}DL��@���qaa%�'���l$���vC��Qk�b"Ŗ����&,��f	�c��:&�ϯ�k��;!�ג��yD;��[.k=2���)�n�o������~�TT-�ϥ����α~�b�ڋ�`�t�פoi6	Eg��r�[W:b�M�ƵQ�^�*�C��@�Շ��A�}�R��ĕq�feJF��5̟~_���ڝ㞑e��a.B�B��-N7�ҹ��1g����P�(y�f#�q�J�'��W]���/9�@1ᶈo@R"������M�;8��<E��M/l�����w����L�W��q��N�1���⦓l$�J���K��@��" �R������s�bu(Fi����������[I��T}�AD�G}=t��%8�t�P���	�I���~�Mi�	��1�����z�>��BÛ��%S��=̀��Ĕh�c!��:�%At�/ϕ�r��";����l�E4[^��I�.���raix��o�@z$���-�@_X;�8QKeqM��/�0��06��Uh���"��s �;'��Y͘Fx����
E\��Z+Y~��'"�	�{Q0D�.4�`Q���xw������i9tb�Ĕױ0Q'�\˲ݺ9?�ɞN9�b��S����x��@��	rS��fy���|~�6�{^��~�3�J�\���	F	y,���{�p��A��UI+��MY\��]�ռ����Y�2_���h!���y��hsz0A��3����$I�qYe���8�i����{p�L�V߿6'�r���kvx*be�^�f|��TzH���g�������0��-��P�t�7�N��ԋ��d�O���:?�1Ӣ3��$Sd�AH�Y����S�d�H�nisbz?Y5qC�	] r�k[����W��.L��=�h���Զ`��'��E�������3z��4��hzuY��S���@x��amR�஽��#ز!�r���w��0�,P\��wFQϘ!_������0|H��˦4L��ky0Ӵ�=����N���IVy˗�B��?�ݎ������eRl��<�ӌp���=�U
���	�(��-��s0Si��������)�q~���������3�2��V�l��x}i�ٰ �ӧฌ����y�Q�s����(қ�ǵ�DoOY�;�<4�ݏ����0�m���t���5d�ً�N��@4`��7�M�H�z���Oqܟ��Z̤�r�MW9W�Ѽg=]�â��d��4\p8b��Z��v8 �9�Sa-��Hq��	���ծzr���!e�AG���}��f���i�f�񤩖4k��½�Vӈ��V�\&m�M��.�����V�X��b�����1?�k7y����jؤdt�@�Y63��uɿ=�Ȁ�=�у-��CƧF�o��p���)��	��:�dl�w���	B�W�%�qc�?�m#���3��F���n�lU:��}m_��� � &����pH�@�K�x�VN�`�hD���^e�VT��v����x:AD�Iy]ǿy H%�3	�f�t Tt�-^ͷ��*��{��"@#|��Ve�	B�V��e���.��� }��6Ծ4rCj(�k���#\��׆Y�5Uٖ�L�'r��Ф���-ۘ�:����&�B����r��A���`��caY��Eջ<��Z�ƝE(���ؕ1�.�!��Z�Z���e-��Z���V�rg�~�H5u��\{֎~9��m�~\	-ez�A�\5���\j���\�/dă㛥�x�EcWZ،��$�gi�V��5�N/��;�R�t�ʹ��jz�i�KAx�e�@���C/�}�ʏ))-{����zCp�����}1,(��~�����NAr���E��v�G�lu�� �8��4
��X�%�_E���GN�GdK�)�ȱi�\������6@`_���_�g/88�_���N0�q,�r9�@ZXa��\��F�h	�rP�H��tU�L
��T%#}32/ 1�`q^����=��X�z�ʻ{tT�d�8�P�t7��>�;8�M��W��[��� 󾳩�ԧ������{㖗�|_U
yl�r~P�,(.�LYؗ����	�5�F$G@�(,s���#�	1��(���%=��$&��2������7��-!�2F.�r�_�����A�-��(��r��[�~�ܢf�I��c�ֳ��_3�֊#X�V��Dt����'��0iL���f���ԫ��	zz��/�m��^�,��-�	s�F�����/��Yi��S��Y%�e��� �E�*�!����bJ��W�1��kx�n��0���S٧a6����k�%��Sm� ���Kp+��OA�6̜����uy{"iBE�/_oJ�ݱ�� ��>���PΣ���"S���7��6]�[�_�3b�����B2֟V�"|h�5�wc���Gv���{9�f}��ӥ��*q�)~����&]�Yt�w�T�m��.i��~n��|q��vm���X�$Ŋ���T�D��)�k[ߥ��ivq~IkI��]��Σ�l�hC+�|����:���~*U������\�^ܞ�4��c�1�w��J��0�q��P�j�X�Naxw��@���d��4�������겕d�ՙ�z�L�Wʒ�VR�[�%�VY�T��i�z�Zk��t�����%ϛXŬc���G��
�0,>�B�|,�f�!�::�R�
�,���u�+��_������	ɿo,�{`=90Toa��6����x�6��U1Ȋrͩ���nZ4��8�]cgCH��尿����X]*\�3�$�z������m�*��Y�g`�0F��
w/;b0:'��n�yLň��	�����%D���[VsL���� �J�3lԙ�P��ؽ��ʡ3<Y����D�\)�  ��������:�j��!g=y��o��,i.���h��Ɓ,�)���U�^ֲЀ���g�!]//1�s��ȧ���KiH& � Nٓ����\���O�1����ߤ�ֹ�����T#���O]hQ�GlGJM�
I���g��[V}d��}On������<՜ K�G��pګ�����R:���7g��aa\h������Љè�ȓы��ȟO��^|�7p��տiJnHu���*�k�#
�R���F�Lh/�i|��F�v��^���d�v�Z�:7.Z��c�Q�K#�<�ҟ^�dS�}�9�K��(��^)ަU�5=$����ZQ��n���̥u3=��z�'�Lf�ɀH{�>�A{S2�IUN�6�?�OO�#�J[Ǳd��C�����lC�ҿ(A�o��[UV���H5A����+S͗���߬h�(&8<�{�R��Pѱu��wjg9��H����Qa����R�m[��Q+?�cZ��eoum<8�<�1(-^{X�3sJO����K��ʮTC^=.F���d5��&�P��K�N��k�u��	��=��"U��(?�L�6��Z+t����ѐ��JlBA5���:��QK.)������M�}*Ud��φM�jf�A�^�o����$.�K���m��?�1r�ڳKZ����^i�&x���Q�u᯸�SdضUq&��?��L"�k��#5\��]eޒg��;�i �Ղɨ�S���2����u�!ma�4ޥ�"iѠ�g�� ��L�I�C-C�-s�̫rs$� G�C>�u����oҰŔI����R5�Xxȯ;��Uo����+��Ɍ�K��؄�����V�|<���z�s{��'�i�<����Q�]��(7:8z��8f3�n����r6g+΢��DW
z'�l��jOR�<�P{��]��>~gd��]>/`Y���=쨸G�ZEebhƎ֜\l�T���=��k����9N�JP�U�!�Jc����y2Z��4s{\D��R�����Z�q.��zc� .ě,Y��r�������7�N�`m�H�?����6[�0K��2�,O��!��^�ZٝT��hqF,�!��K��-H��!��xS��ů��+����c$��D��MjQK��+���Og��8�Z��l4�h�Ǽ|���Y�R��u\="]|γ/>}b��k��qiӓ�`�p�q^��xj���z&ʢ�}u���K��.����0|d���2����Y�D��}p���5(�)g����ߚW���J��� e�»�ڤw~:J��RZ���,�7��5cL].�t櫧��)4���\r�i}�$����gr�i�9�e��;>� ��Oc�����Դ�v�lr{s�!�(��೥���W���\����_v�P��Aq&Wn(ą\��r�;���
�:�����oPu���?}b��T��s�h����㩟ڐ����dp8��eQ�|x|fx��lf��|���m��ԙm4��Տ'�&װ��0C�� ��#�V)���U<�]�h����W�K�g�8_�׏�Ư��������0@5�HN����/�`���+J͘e�-����(�>|"G:@��S`�a�}t^N�L�WA9�R�K�[,.���l�H���0���*���l��1�?B��Fs^`0�K��(�i?Ԃ]�t���_u��$�@���&��srx�O�/����aQ�q��q���|Q�'+�@!����/2�)c-�qg�;־�*B�K��ӛ~^{Py~�5�Id��]�|�����û�\%�|Ƞ�Gax"����=
U���;���eW	`m��+ؿC]]JV3�iB��A�5\�s8P���J�UwU�C=E�U� �8��7��8<~�Ѫ�Z��9�o�5g���>�^z�[p�j�L���a�BY�t4����e��K_-.�>Ә�F(i|(� m�����D�Ovl]���d4!����o$>6�]��,�a��'l�:�;�mPO5��F6�"���'hJ�uּ_��څ�mJ�{PՑ�B�і�{NU�Z��F�}K���9p�8�TFcRyJ(� ���i�B���#��?��1O�X�"�!��Rjg2o�3W��<oy�~�oBHsZѯ:���v���t���J�~�8���VF���Ii���5�����R��CB:� aF�
���*���%v�*�Mx�������R� �~�3���*��C�29=��>�)2r����3K�"��Z����yv�� C @�U�b�'[r�?/z��0V�DQ�=�e1�_�f���-�Z�ˬ~�0j6����sXm�"K乂�Y��L���ى>uF�ȹ���n�>��۾���.�o\*��Az)��wg?i���*�$W�����k!:�?E�| ��E�� �;��;�`��4M�J��'̐��	�5$�>u�T%����jse��>ޕⳀ��h�U5n<D么_���Ы)�~@FFJ��c~�>�b$�C��`�?���G��~���Ĵ7[�L�C���L���/����e8aQ��c?�՟�
/)1P�e�D�9P��Q6(�(�hod�gǞ�B�VTW��P����u�V�U_�ʯ-�J���F�ŅR_�	���
����߅M���>�?;�-6�)�]%�� {�%����r5a�2�Lp��ߣ`��:!��9˓��wn����Z��^ᕁ���K
��x�Q�RA�D�;��3�}���75� �����������vP�M��!�[@蝾�x�������<ĩꍐ~'0�3O��B�ۉ.���ѫ�$�~����揂�yF`*<��V�J^�IҎ�&���KS!T��jՙ�2T���m����wGu��Qa����q벶»�^������[���"y�
 '_bh������L_�+6佴�����7���?ح��#�9	���I�6d�(��sN ��<g���A��-�_gz9X'�^���v�S�F��J��!��9��V�+Һ����6�� �-�m��2�
��K�su���0r�{� �OB�̠���G>*�ߗI����tX�{9 ��2�2�}%���>�I`���A����@�G����M��v�Q={%����Dk��#SL�?yo��8v\�U%��8�l�5�X�����mN�S���M_2yC�,��xA\|R�o���b��j��T�������m�oq��B����n�Š�׿�V�s�D�fzh��X��N�^�S5�W��~ڑFv�p�k�Io���c��<M
^�mF�>�m;|+)
��Te�ј���|A�F�O�b��7Zٞ#yWUY�21�H��ڬ��|*A��_���=},�����\{�,*�C�����Z���K}�բ��\5����C�*�ҝ���`� ���zr±�^"�'�2����{�l���O9��Y����R3nT�P�9q3�	G�)9ŚU2gb.�`�bw��>� ��j�	�:.���������E�b����HN������ō�Ӭ�Z���߅i����b �Z�k}�/䣳D�=]�S��(����Mg���m��p�I�Y� �xfԍ�(�ҋc�]����.ml=R��bZ����z#��Sp�u"p�K{��8�uS� ��2���T���*����W��1��*sA�(�|��X�j��2�s 4G̸���qk�2a�Y�a�������������P"΢�Y7��M|�Y�8Y�����w����-k$:&�$��m��j�A��v�,��UK�D����a�AvT��G��
�#1��!ʵ�i���[�0����հԅ������7�U�Y�m��-ך��,3�ɶ݈��Hl4��]!�+8{�NG	�&���ҏ_�Mp9+�؜����h��eWb?��}T(��ě���+�񜂩24����eF�4�������'�\WDq*lc�z+7�C2��3K�<�����c)}yDg��b5�i��y�,Q��� ���Ej~�L�BЌ�d�y�Ed̨�Fg��!���H#rg6;G��l� ?�C��-�̱'k�{���C	&ˢ���7�r��f�~��-o�⅑y������3?�PdYD�Y&,/m��Tlbi ~�Ƨ�nڛű��ne�3(���dT�)��|M���H��ɓB�m=&��f�}�RO ��<��Ѹn�v�8� �PZ��p6s�NrJthP�Gp��	�x��ǔ�EUDt)�:q��HHz�,���#��j��b�q�����t�3�":�b�2��i�����Ņ�� u�>oY���RH�����8b���9il�#xQ`��ԧ�ߖe��zy��F�#���dwn�T���'I9n2��Ti�k�[��N�P;ƣW����p�@�"��}� L��-K/�Ц�r���F�N�4.,!��+����;��	��t�Hʴu*A�^2
���'�h�W�\èe3E�:5�܀Tއ��h�/G���j� �mpc6����;W�2(���W��Rݘ���qzCm�~�}�j�C�������K�dn�x�l#iK��ĺZ�(�*˦F��ǩ�]+�c��P��}!�2
���~�#L8'�L4�*W~�1��w�A��멾�`u��A�h�ޣ'2���O��h�ݲ��@)g���XWϖǬ A4���Kz��c
��2p�G6��c���vd9���¯�G\���f�V��$�~TjH휕����r�59�m��,��:�ߗ�0��h����7ӓ�;�7zܭ�}͓���O:��FF!���O3U�Fj�����wi�����I�4P\���D�n��_�i����������J啼 ��a�W+���g\�����rH�T��d����<��t�Ku8�^{�ǹr����_G�W~dI�G���D	���Z�7\~��=����@y��p� LI��Fn�H�;��Kz�/Q�`'{s8J=o�!]W�ܸGH�9�KR��J���"B�@�ř `Л�� ��v�Hg_��<�sA�~`�`�d�R��w,~��|�q��v槎{]�ɼF#���'�xͪ���Ec?!���,>͘N�@'�şx�@��������z+�S�*�� N�9�eS��f��П�:j�搌YmBo)
t�&!�ÏЎҲ���ReJ.�	���I��&���SbK�;<~�St���,2�bE2��<�im��Y���~}S���gnZ��, H���b��z1����z��v����MdÃ�8ގ�j��~�|����V?���ZB
m�t][S!�ݒ�~ g	�,
�Uc/e\<6�޼�fH�[�t���V���;o-�
ۄ��ùR�&=Q�f��d���_m�H��G�a(*�ED������ٝ�Z�b�@��
�3�G-���~D>!���B,����]�I\��
6�۸����������ў>��a���Un�D��`O,�h�(��,#_�^h���,
\��a��������m�!�[|W$���`��R����qY��Tā7�$A�����|J�d�� �Ӥ�a��7�3��Z$�'xF��8�ݠĔ�Z�1�!��7�a3���@�?Z	�F)�}?{>�D�����աi��[-m/�؜l#	:������>3���s������}5Fm^����;+�6���^byOT��a�����U�վ=:�X�	z�;��D��(a��ç%��=p{��g�dYd�����}��S^
�Y{;ic���,���^(���x��(�#�ʆ�|'��ç�����i�p�s3s����}�w��T�a�W:Yag��p<4�&�.������}�/����A.B�P���EL"\���}M�(?*{�� Z�p�Sޱ�7[�1&z�ֲ������>���	ȸ�H,L�����F��1�@�Ά�,0���u{�`��Jz�v<� �j�5�(�D>�Mv�Xl���Q^?��W���a#���,/q O,�����%)�����S&&J���HP��4a�hf��U,o���熶�:����bgɘ�b�  x85a�lt���>�)m���z���XG����f���1AX���C�J�l5��$�m�y�_C����uE�����r=E��q���\7DU
*�T���=#�Q)���ĉq�҄?��=�D�M�b�;���lE_���N"8cy9��d�ůc2I����)�b^y���%lx|.K����4�@���w8��9#����N��Wڤ�R��@$0�mؤ��Sg��H||�����ڏ>���Y&
W�Kb�F;�|**K�15��H!$�6�H�å�p��2Jv���lB�K�JO�������(gAl��r��ЉLz�W#�2(��}�4O�t�����Ů�:��':��v �Kd����1vbh�/���~܂�7���&&���t��]R�H���O#���;m�Q~��UA�^�dh=��l�#����a�h�/+"�,��/�0(�'��0�����՛e�Ƒ��+{�r�HH���U&�-<5�w��\J���nৄ�$�Y�"�W:�8K��3r�~�%��Ὄp^��t����fy��.�gC���'�G�������PhAfܧ1�+
����W�cVrnwq46���B�ep�������ٖ=�oV��	�@�������hpQf`�2�hT�Z���3J����P/2N��`Y0���Y����ǸeK��=Ѫ@|'V�G�������R���7��v�Nh�y�Ѱ�P�TnK�Km�n�W���|�V(�m�%<���Tx����M�yc%��50	��-F��	Ȥ&l㇀H�j�Y|��OQ�$��kU#�4�Z+`�\ TO�c����sy���{-�[0"C����c.|E�\q�(z�0f�(�������Y���;�>`�T�e�c�����s�S=����<m C�!c�0���/h��ഢ2���i�أ�X�
~dr��[��>�x	����?mq���%rc��j�ʒ� �O _���7�f
�b���l ��.D:��G��=���}nx�����y�� a:P��u�P9��i�rvn��#3ך��v�t�!c���@�`��oY%�51PU�R�陣�L�w�t@&'v�MP�m[N���@T>��-y(��u�;��n|5��@hH
f0�3ER%Z҈&:�A��ii��Պ�m����-���d��J���������g�$��L#�+<C�:��T*v�$���J����P��R~z��7�K�j��~���J�$Y��*�ihY]m3~B���h�=I��:���n%������$�K �I4Ϳu�7^�4�:u_��h2�L��&l8+� w�3�x�w]\�j�s����'�ղ<K�ʨ�)�wZm���Z$��K>Ԁ�
2Q�>�H�}eq��)��R�7�wHgi���C�̘� �o@�)2��{Ƞr��x:��(R��X^r}��L��UY��/Z���=?����|�&�D�w���V&<,��9�|������G�?D����k�Y�Ϗz���Z
��;��b��'��J>E�mj [!�&Ok�U�d���/���K�J��cb>f̳=b�&BJ�I�Q"����]G4�v��}~��԰7\���!����%'}��R2�)�N�6}���B����a'K/.�Q�a�XY1m{ �����]ñ�"�������3T�3�ʙ#Xcn|��g�~�@�R����h�8{`w�Ce5N��;�.��j����<]O���]�c� �*�7%�K��¯�-���cYÓ���ý�L��b���	ػ����/e(�g�J9<���笣�̆�܂Ow9���A���<M�b=e[o����?z�n@k*E���H�_K�T$���#���rL���k[�C85W�%[�STu�/5x�=�����[F(J8���8����V�V�ԭ4g_�tB��kcb�W�H��X��A�T��Y�W�t�#�S�KB��m�+�2��M�$E]q�7�\q��xPi�+�"IGG� �S��K0w�T�ǿ̊뚽��ѿ�����1��8�k�O��uS��z���2���T����R���6Ҫ-�W[�HS�����{����cM��D]e�r�>�^�b22d�@mĉA֌"	%ػ������W;��i���0�3��z�	��෯�h�C��K��K�G�g 6/w����	�͗�f�+,��C�����`��F��.hx����<�v?���~YɊ�{�ɳ镻����zW̷>��f�������Ju�d��U��	�ː�!֭��Ct��U�sY��kn`��Z�;�q�ե8�aYL�zտ���ѯ�«��Y�(����-d�ߺ2�J�D'�gdm��\�!V�/Ԥ��f�n!�5i5����~|�k2��ܿB]>��-��Q�h�#�]X6�J�q/���=�=��o�g����J`]D�Ue�ҫ���sD���SҔ̝�Q1/\� �v�AX��İ�i�o�1���úۡ����(�����l;2��Q��b{�/}�S�P��?&+���BAȴ��K��[@�������̅3��S�K�<t��S�ϡPRM��egڱ������*�V����Y�?�Mk��;�fm�DZ~����8[�x�_��с�?�����Ө�/�/4�����d/bB��c������@{S>�'a�Ժ�P�ᔩ:m�]ի�G�	��!�ZJ��)����͐�Z�e��uO�?���N�>vf�.��1��a��
���G�R�9��.�uK�"�=	�`��\�]�pj�d�IW����:*���©�+��܋���ݰ�.�&U�,κ���;���t�`!�5�X{j��2�W�>.TB����.5�nI�����f
�bѨZpp� um�I�=��W��iQ�v�V��˞��Ap��PϵG���J�5�h���D"K;���f����x�*��%R�����~��m�
��z��ϱ�A�gk�0�u�xPᷯ�n�\�(�*װ�}������ԟڳ�v�f�Ց�ge��v�o�)�&�$HI;��M�Q��9�x�k�iK� 7b��*Կ���eoߞv�:]�C�I�O�w^[���6���#D��*T#�I┰��).��Php�>:�����VB}\����tz�Vt�bEc�_f��wU��ѦRF����B�l�N�i�m�n��z�ҤF'O՝5fO�{J��j���e�aJ�I�BD?�i�¸��Ή��K��W�on�������C���n"!��/�����Y�DC�Y����aO�?���J�x���5�ށ�rU��̠��ԅ���u�:¦�� >�{,���q�bM1i#��t�j��0PpҠ��-X+���>�< W�C!$�����⛙��]�@�-�N�:�3Tm�|ы�����d�BQ�G��BxKL�)=��談��R���TDUo�Q���c����#�c�Y��xO��E֙�}����l�/������g/�a�4��NИ���Uf!��H�m$�W�t~r�59ȏ�`���Ӎ1�bDLqM�QlI���@G$�ȩ"���7�RIu���OO��~9�h�~<`���e#B���)��3 X�l�?���.}��S�0ODk����=�$'S9��&}b��!Z_g�ֺ� �w?��+��[>2�v,��3�iR��n��(�O⎿�z4�!*d!g�l! w�t7�#�ta�a��s���	|�U���"6B��5���PVx
���G#�Z��J\5s6-�I?B��(�7��9/��x��?V��qT[�f��5��~6A���*a(yE�C��%��>Q�/5^� 9"�(`���g>C���/E���z�tB��=�ڼ����A�@5sW�
�r��"�OQda
g�rIZa�bO
Q~��Jߝ��,��ŗ%� '!���MC���
G��� /.2:N��ړG%�J��	�����V�(��ǉ�_W �[w�:���{�Q�{����LY_S�@�3[�#0���̳<^���J�8�O�����K�1h��,�HFc�W�nWg+���}"^?ork���H �����~h��ߥP!ߢ��A��̀�S��S������3������~��v���d�$� �Kd����7Z;���kV�ۦk_n\�C[���ۇS��{|��u	>����\kAY�c"�D���|U��Hֺ�ү�ٜ�}W�B㮴���G�n�uR@�M���� ������,H�C�֋��)g����u?�ߴ�@�.\^��z����s�]���;G��"eH:*��e�� ����i�����X���.�.ǱA���x��c��EP"�۝�ݺ��#Ve��7�L������q�G��og�g�ڗ��B�Z��=3.�_Q�j�����ه'>�[�x/*���{�'y��'���j�h5MC:��Bӧ�@k������͢ﱟ���&t
$�C2w�	���~���H�����{��BU���xϱuR9�@�I|��'Qa�ϙ�yCE��`�wm
��❻L����оD6H�D&r&���bqӤ �3E]1�m2�2��\���<��`���x�5!�<�gxoG�&���0I��.���\=���{t`ܬ.ea&����n�9J�kc�K�ı%f2�7|h�N^1����1��"N�P�O���	o��1r+�	�}��$!{�6-W����S��R6�AKV,R&�=�����Z9M/�WAyPU�Y�Q�=��rX��w>��)M*�)Cy��u�Ij�J=�#ka-����Ê(LV(���5�C\}8��p�E����k��A���֚�X��o���a��{'p��Rp �(�l�2Ì�~��H��¯����:'NಡQ�_rΏ��e�Y=m��?Q�u\�lX�������p�.u��Wޜ��(�H�D����S��Q�.��]>DU�R��������'��[��U�$)��������zE۽~=jJj�����JrRZ���BbG����Q�����Fut��x�,8�ޔ�	�v��=��C� ����h;Ň0�M/��դ��y:��m�;��_�E[y*�Ω�ۡX�5z���c����8��h���Iɋ򩡮���~���4�Cb�&��@�2�c5E�8�uN�\��ą2gEG`LdK���.##jv��,DX��m�^�c^{������j�e����R	��hSS,Lpp��n#\X`�>�$u�m��^x����0���b�0,��ar&\s �� ���Q�����E���4���_�B�T@��s�U��Cpn���f&L�Jп�l�Ƀ�� �D1z����V��Zg˚'��!l.'~���_����E��P��k��Ƴm�T��?�C:ˇ�Ѻ�n��g�v�;�.eAEv�ܯ-7�z��]Y/��J�RXؔ�AI�����Z�@���'��G ����=����Ih� ��xW�"���R����2*�*D얚~[����t���k�-B6_z�R?]�[��%f�P��b��������X�>s,W�QUw|��X�!f��A��'���e���~m*W���r�PͶn&\�#�c)�>x������v����R%c�|����������
�dȺ�p�yG({(�[h������~8r��G6�ډE�Ȣ�7��.�4Vл�Lu���z�-���<�-X�?8 p������4![��xʐ D<��CK�����5�'MF1��X�����؅�#��r��(�~4���QԨ|�7�q�
�N+g|�!�~m|}Լ{ln��䊟jX�5S�9݌:=Ki:�iB&�u�#��,b���fK| G��"�zn���5��9l��;�T�>\Y��~�">��������2,w�Fy�(6������������tq<�>ab�S�e�$�2���g��e}�b�vʗ(}�G�@v)7FV/f�L16�/�Uk�vu�&@��������Z��$
<3���N�Ssx�(@T���ZG�q�뾚�}F�\ ���nn�s\����h�!�ĶfP5���n�#�4~�G�(Vs[�u���h�g��U-|{(�o,uJ��͇�C%�7+#֬j.D#�&s������Oi�*���[���8��>�LJ��)ӆ(T�8��E��k^?�T�w�Lp�*���&ԁ�L�0i�H\rA~Pza�Se���lA�����z������M��Z!Y���{Q,_�SC�옸�D�k�2���V+q�ߧiL�I���,r��W{�շ�e����)<4<��F7�nZ��E�����si��@��:{K�=�]��`�FP�� �݇$e>	�gj�F�yW6��ri�D�S�C�E
��.9O[�/s�b�PIE�<y*�`�=�q����_�:�&L��З��)�����^A8�yѡ��$�~���W,��q���S�ϊXOk��_pL�����rR�(��7Z�m��Ն�|Q������|'Q�����x�"�\ud@�[!��y딝v/x����b[ Dh�,�#���w�����{�)�t�Z�O!�nMs��@�B'���]}"��)�/��oD��,(�dI!�Tҧ����R�flT-O���=UH.H""{������_Z*3˱i���_��P�~������eg�ZkD�����@B����|3�_m*���.fC7�t_>����4ɩz��q���W�g-��0����w31�|�Ajg���f���>R��0��B'�������<�y���/�@d���;5$ז^p�=�V�W�]��%�7�^��{��mP>�.���AG�yO�x�K���)G��-f��m����ҋ�/����f�"p�����|l�(�]���5�I+Yf��^��B���@���v�@��9,�OY[�UkeI4�y������p�jꕭ?�sB!x�m���v�0�1(�R�6N���B��~���+,iЫ=rE	�J��[���u;`GǎtgZn����?L���ę|w(���a�SH�#��oj���u��u�Gs�t�^(}�Q#�o�xd`	a�41�(���uW���Y��]?F�9B=8&�.Ny�%
H�wy�W5LG��a�#���(�џ3\y�F����L�X;����� �d����K���[�����90�}v5�F<E�#�#��=}vQd�:�>�>LJ�U���a�_��-��Z� 6�0�	N@�c�AN��3-��p&�z�r�p�y\+��j#��kw�'O^1<wƊ^�G�沎��^��ӵp�x|>@3w�gb��җC�5��܍�d�93_Wg�v:I�,ٞ�	{=����8�$�r������i�O�̟�cڹ�ك���&�Q%3I����fF!z�
�ߵ�K��t��&�P�9�]+Y��P8��<r}�����$�N]?9�r�@a�=V���PC��8p>������H���l�<_��]�E�|�.	m���و�_֕�]W���s��_!(dA����K�\���+	��ʣOM�}� N��OU�L����&!����#zc���ҾO��heiެ�]�3�^g���.
�����/M9_�G�ɚ���T�S��Z�wL�{\2_��bC(I�%�j�U.�"��u2n��Ƙ�b�+I꩹?��y��
��	�3.,k�-�C�e�]����g`���K����R�T�r��7TL��/�@�_��4Lq�{�
�·jXJ���ſ�;d�vO,Q��6'�̖*�O�����^n40 ��o9*Y��5>0��H�!��	s�*�ws���?�MVh:ߜ�����ԉ����B�b2�5s���+-���e/3�q��{b[���9��Q���Y����f.����DU=:�j���"��J��ɒ�w�5��Y��k`R�F:�ݎ�gs �/4h�!�*�> V��_2���&i������
��z�0�L�Ɏ.�~�K�B:��2�j��i�.��Z�եO���]��Y�����X��Ί'�v򨆞�� �ೡJ8b�P�\<4 �/ju(M�w�SU#&k͘�c$ꬶ�����Ly�������4���X+M���Э?�YX��'���U��N������YO2���A+�U[V�!���7��c�)�IY��(�����_����C�y�ɌѦ�zz����uf�q̘H��~�*kG�ә����� rO&"�*y��b�wOa�/����J�v��\���n�ڟOM���6P*tb��~m�[��L���1�r��{pK��_6����(����b�[��ae�4d�c�K.|��A���$��F#�g�]�~�M��F� G��?��kp�f�c����r(r��c`��hʒ�7(eoĭy& ���jں���T�q:ۑ�~�Q����0���?54��2�A�x��W�����-�+b�,o�꜋��9�v'��Q�ٱ_{��i)Ү}:-zmo*ˊV�|X\%VZ�����G��Y��!��\a��H�A*��Y����k�26�S-�B�E�UPؖ�m	�)���OH1o����%����@^�S6Ì�4�bw�	5�T�=��^�`XlR���c9��"S���&j6?8"h�$�p ��u�l�3L��O�Ee�+$�q�	��mb�!�)�4�n2� �⒎d���k`a�<zd>_�
��-���14�x�n����X���8�jǊ�lc�(���oMW�����!�7�Q]�."ȃ�0�r�<�7@�-ґ|���9dOF[��'ѝ��(�Ė�d�|�pX�-WF�V��s�ښ���9L	�`9. ��%�����yd�@��{�>�&�{�B���R�2Q��ZM�ލ�]�E2���g�"�f��˶Sp�(�!��,��	��P�D?
ZL��{%����H��%����N�b�$�'�y�����f��xeW���I9~���P�':�H�(G�=��H�&e5�M/�;���Mj�CJ�!��Y&}��d��EiQ8��-9�<cٱ��������</q�E�fq�N	S
7���޾g��j�4ãh�/qJ�g���mCA��4$�Y0N�cn���ǀ[Ѧ���ꭊ�԰�*"�ַ���E���b"�Vm ��A����e��@ޚ���ZٮvD�^��MT���Z\����b��cC�i��#����uj���J���f~�� Ӓ��b@�
�����9��Q�'������4v̍�ĤF' ] ���t3wÄ7[�p��vGv�ț���ޥl%%���m�lX�J$� �N'��<�^���%���	�IӲ�	���_:8�|l���"3�
?��>�U�Iݴu�ѥK�X�V�d6e��*_#�3��"���Iu��(���?bu���p�()|��?bΗ�X����9���<=뾹����Y6��F�&Jw��r�f?`0A+���d�����<MU�B�QZ� 0 ��c��J�ۇ�pp$�x5#����c����I��=�x��4Ks�&�{{��'�
���ԉ��U�B=��_���W�%�5g��K�|,{������s������Hg��A)��%_N��%^�H��p������3�/�l����hd�R��y��)�;I:T"d}o	<��)����bgCp�)N1���FJW�$4��2?�ϳ����׎�J��X�a@&y�Y����A��,]go�L��:n�i{�a9�bx¸4���>�2F("b��,ȝ9��6�o�:�����EZ�a����@�*�j�)]����.�B���C��@Sr3�x�)
٬���م�����i�=a���"YK�оG��:g��O�*�X��gUv���&��x���
�����B�fW�R�VP��_��+Y�&K�X�W��������?����M����5S�ɍ�A"薚{���7����@�@+ח�
`ޔ J6�$���A��$�Yhx��f�i~�"c��������w�ݐ��Y����X���aE@s�B���J�N#������2�hDm�L�
������o�T���u�˧
tT� �Un�G����L�OS�����Z4R�͜�~�em��h���ddP�(�	�bV!/ϒ����&�b��^U���V2��Ȅ���@]\��Tp+�m�g��
������F-~p?�Pg`ߤ�Z��0��u���3���,�kz�@>����ĸ� +����V��/$�F��~���/n��M���x�����Fw���ƶ~�O�$ֹx�_������Wd�� ��@<7-ڼT^.�	+�/�,�g�A�"x
�S���0i2A?�ZB�ӻO9�\ğ�*,?42���1�5Px���R����S����C@�m�XM3���I�@��V�8��6ݻ}e`�{�9恃�f��U�n �uu����{z2ۘF��{d�V��>`��������o~����!B \��P�0�)[���͟
��eTE�[��L���Su�;�KGE�:����+��2��Ĥz��H��6�.1`��H��ss��L%����&��Q
����@�5w����A��٥P��c-��oTt&|Z1��Z�4���Wx�Uc�t4gʆ~l�2�a�vk���_���.`�@K7�T],��\�1:G�Q�gt{�ĲI�7�2H�Y&��m�t	h@1�
�Q�|2�ݴ���q�*➡��qк�@%�#���B���A�X5���գ��r���E�����;ŧ���bj�y�a�Q�G*��1`�),ka�tO�|�[[đKO�k��Y�ku��J )g�؏�}�j𪑜Z���%�ϛf'��� ��ٞ�-���/�E���]�X�ێ��3--Du�4��G�����g<�
v�
�]��L,)�Dv�= ��۟�T�vګ��!��hw��M��ht�����`�h�� �B�/��[�v�Q&���o�9&�03�
_��j�X��mֶ�J��R�Uۢhg���$+��M�#������2r�	���^hr��
K�{}\ȯ|���6e
͌I�}5�suR���q�r���da��7�p/<����giI�e��(:��,k���F0��2+'>p�Vm�,���F� c�Yl�By�h����3;-Ǉe�7t��Ɇ��*�Gբ�=�Ϊ���6�(9~;���:�Y̮��i���'W�M�)Y����
�(W������7꠬r��H��Z�@�;�wf_��IU�G���Wݜ���k���gU�w<�#D{�O�Er�v�
�G�b�S��鮪THDni����Ӂ�-*b�h�����U82 8f �~���/���]ӆ���	̴o�ZÑ��P�y*p�����)��)C�q�Zz����ҏ,���WT�����V[��u^�����Q5@�L�����Lb��(at���8�#g��4���K5���Y�d����H<ձ��{�Q��kK���b��ZRǭ�����W�[{J�P"]�����o>���m�s��P���S��<k?����H�M����Z�`�g�F)�w�8�ʮ�|��51��6
+��ω� 8��池\D�~FI��9��n��&E/Y���u�)�J�ч۵vg�P|����)��?k�;"u���]���h�[�Խ8j�\;������́]�s��7?����oNqv`u�&�~;�=�Ț5�-��`\��)���R�&��
��uY���^����7{��]��w4�ơ?��uU��d��a9#�$��j����B<��P]�������A_8�L
�a���t��FR�.Ѻ�q�I��Q�R�Ju֒m�=%j( �]y�b�U��x�S.�i���uN��V������h[)_K�pt�����1���i��[eܗl�Aty\x�ank�D��9��{�ջY�h�>}��Lp��q��pD�Ex�'!������xJO��EHgC��9ozK����5�,��*,ޤό�C+��7B�]v�i�X�D����k��Y�,��EYq�(9�J>]Q��,��5,��C롎�����/c��.��]}��f6�H�ۦ/��p� 	׃�Yf����&�ܪ! ���2���>��.n�v���t�,y�%��&Mo&�b�C���/**VHjI��l(��"秶vȫ�U�}�K�C�k��E}+�"��h��]��p�:����:���	�(�Cq�]+�p�p`Ρ�6K��B�^�zu������L%��d�������0��ba�((7�5S�Y�{��_�t��8��:A,k.��*|]�<q�N���
��<�Q}�z�%7�/��)��vHc�#p\��vE� �N�c|Xj�����q"����.���g@�)���f�N�G�Z}���A��
a��M�6s�����8?}b�0�N`ֲ�����/�8C��R^��:��r�'�Ķ֓ne��j�[�+~_�j��[�Ӧ�N�����r���OP�;�*����X�=|��]���뢊.�
�\��d��J�E7+����Dt�ڟ�;$���4@�ۨ��p����4��u
K;+��4�-u�޺U̺�pÓd[�)�yx��2E�]^a+e��q�8�1��S�����P#��Ⰿ��YV�T�:�Y��t����Y3�Cp?�{��ܑ��¡�cf[��_��5>�i���ء 