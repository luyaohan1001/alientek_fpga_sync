��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�^͉�������A�������H�&��&��p|[��zpDI{,E+	Bb|�w��b�Jq�J�ȇ���4����������/��})I�N/	^�`�g��p�|�O;��~��7+�[�@�M����0�ѯgʹ��j�O���נ��8��]��XV���cCt\u�+�l�/��[\��h ���pw�D�{H�ί����Lt�Υ=¥(�W��.��a޵q�����o�lQ:��\�>u��w`����������ǽ's�B��&Wn������R���jµ�7��*}$�e�-�h`��m�}\�T_��n���~I`�sVζCyts����x� ��آ9q��#����H�����K �W�͝�t�Դ=sC�j����x��E����P�,<B��"���	��餈�K���=RNn^ۭ�L�ʢ � ��[)7����ATKæ@�q��E@��T��h�8\�XjRPY��ɗ�	�?S�fc�[���w��
�n�-�լ��2N'����O��Fr``���7"#rj�ъ�zR-�6����]P�P��FYs1�
�d������[�?��< /e��/ћ�G0���N��=r��\ƍP�s@��#S>�����R������D��~$��b��B?��T�Ô�+�,f{���(.�������+��ch�֖!E���Dn� �; ��5��������Jq<f���^Mz)���-W5������ۣ,�K�ч�JK��g �����?jt�:6���"���G��2��:���G�/M�Y����\Q���J�����6`�A�4�5�Y���S�{���?o�b|W�Ԑ�5���(SB5e�A���!��L����9DM�$�|�
������5��������:/��_4�X�0��X�N·Y�О�j)�Lec=Z�ӓ޻P8��ć�s�����	I��l*��曏��}�r}��>�v&�@v���n��yA"ׅN�^%&�m���@"8/�?�,�_$Q��:��i���	��]N��P=ԃ"g��~f\,�K�s<�72`Hp6�1��{��т�����=�kG7���u�f��΅vjB��u_���H|�E������F�/�3���,��
���b� �� ff;�`8��gd�\u��7��1#��(K��W*'�H�^�+p�tk�Ώ�����N/&Yni`ܡ?�>$���IX�qP�Xy��fH�������p������5#��k��(� ҝ�͏�|��W_��y��YG�~�JQ-�����-�=Y�3٥Ǿ�.�%cx� ��^ �K��A�������U找O��>�g̀�;<C����iy�n��4Y���a��'���\�J����^Q�ўa���p2�e�L�Cb��W�M��m�����R�3�c�z�g��k���K��y�oY��i�p�/�*¸ %ԣ���d���zG�|��
Q>��E����'е�8OM���`���8���IK�_�h��{q�0Ra��2:?ی�?a��#����m� �f���a���8C�3������+���q��F=��`�eK�c�i��� ]�,�]t�@%� �$o����5d�[|�\�(�\V68��Q2A!���խ�B坞ٖ��w���uCC��,��"	z��������4+�E���W�4�^_��E����ѩQ�����7A��yy�
GQ]�^�Rա/���xk%?���}l�����.'�X�t�q9���4��{H�/�Q�_�:($9Il���{��]6pZ�c^�E�Jb$�� x���aEj>��~��yޚi�O�4��
2����P�hq�[F���!���K}9ў N<�-���(A��?�=Ģ��#�z�:ѻ)����c �~�r,dTZqc�dX���<(<O;_cJ�k�f/�Y�f#�洇C{Jt�3�8�:}Q8�jt`�Hy���8��h.�Y���[�s%؀(�N��LE���.=�fڼ�aD��d��)��?)C]�˻�¶x(�+v�"�_G�/罗S��d�\|���Ff^i����H�r���w��t-��&�+��G9G6� ,����s�H�)����rW���ʴXr�A���*粆��������9�W-��+j-�D]m�FIB�I������z��Af/�����$E�>���Z��Ѹ�o�W�^��K<�#Z!2��f�Y�������E/`O5�ҢֹP����������a�w&��K~a��N '�����Hi~��R�a;�s �l�J�j��/�e|�)��w�ks<��g���!��{q���cBE�{�+EU
F_>�%���{���k�錎�E�z��Oi��P��"HDy�4� $d"���f,ް� ��n`��X�6Ĳe��+��*�
y� ͤ��h���ec�'%�'�-������*R ������i��:��+��T�'�4�J~�Z.g�}�֠!�k�_ 0���(���!�('����B�����oC\��=��� ��x��[͈�)Q(�	N|ՒcpC�f	����lsΕU��os#&'��'�9�6���1&��/�m�T3�d��� �B_��;�@�*��$w��S���������M�jr��+K5����l�J�D����ۧtc9�!=C�LR���"�l�h=�ͥ��Ĕ����n�5v�����(2�֭b8F"���[�����H��[l������Jq"S��w)t	8F�����cS!��R<�+Z��F��;,�]���{������P��!>�$�����������g�i<��G=�X��8�����<�>�!v�'�u�a���I��zǘ�|��9lJh�y���U~Z���p>�Cm�,%�$�ן;g��-�1�<h��"�NmVО@1u��6�fH�~B's+kB"�z����5�p��
HQ�prqq�#�)��*6�V�1����KYQ�Қ�}�[���[V�vĕ9�37KW��_��75އn�EO���c qG��
��h˰������c��ֱ!�dZ���hB*��u��("j7��M��t���mi�'��)�
���97�$r�a;%]�\w@���7m�Of
-sC��Oh6M�l�r������v�wo�9G��A��?��T�bګ)K�~�����F��Ά�;��V"��0�G3.--��<�!�R.�����Sl�5%��%�Z<SaT.g����/#�4ޠ��\��֊��S��j�ur!Up��- !Y \�2)6v�dW+���l��)	����H������(���W�l�3���0��:��{��.p`	���C�HR������0�R}tӃ�|j�^��a�ḧ́�f�x��گ���䕙vmT��Ib��R�uV\��B �%x���G�=�[�}�q�l�`�)��.qU���"q�����7c�{�1�D�p�V�e���ԯ��s8�n+q��.��:��!r�Y���Ⱦe���ū�����޳����Ҡ�I6���C����$�H�h�\8�,��ֳ�u�+׼(aA:e���§��AV�5�qx�SB�nF�V�<��'���k�1��I�p���j���A���i�$����evQ���G+	��4��������]�Z��M�z��-�ѽ>�����H�/e���
�_��i��)J�<���̐P����6���$z_�	�H%���r��ޣ��]xx�(��QT1����g$�U�I������%U&�~�3J@���;�_���l�P�a{�B yE7S[��Gh�r�e-��֔S���}[��ƌ+h�+��?��)-�
�2�D+�Ћ��mO�Έ��Bf:]���å$���G����;�r�bl�$�n�㦯����Ss�)8�;��-��9:U�JB��s�sݞaI;NëB32�_L�@g��R���Q��k�����rZ�u��7�?gǐ"�q��*����K�����1L��Ie�A�2H�]8P�ȂӒhNG���T�7����"v�ލ>u+��z�P�>/�
�@�f�g��x���y�@�dVZ���ҒW|����u�o�����
y$.���V[����dk�v#A:�ﬨ�2��Ek6^��+s���|t1(��iXi�`�3ф&.39+�@��u���H�B���r���gLn�������SnKu��~�.���6ۻ�(����#�!�'���Q�Ι�o���4�I�$���r�̾��qq��w���Ŀt��K&�Gx��#�8����ė&�V��(9�yR���<9v:�x���F�V��	�'���ҔQ����'p@T�u!e-	��k���:��~�����
��]��x��UA��c�g��]���!�-��40�������Vf�ϓx������'�{�.��c�}�%9��Łԡ���lٰ���-@�D\n�!%1���F��$4Tu"]8/Z-L<�z�n~����N�b�)	F����uiF��2)40ĵ�s\FV�:L��y�!?ț�Ѵ�L���Lچ�zqM��N���B�	��}��lN���1F�Q\��-��yr����@�!(gӌ6ei���G]���6ʘ��Q�&������1���U?�E��k�CV��A;��!Z�7���}''k���P��t2�1��G���K9$����m[��({�M�������+����~��T>"G䙎�aK΢�^f#�g~*L��bԄ_.�̥�n1-�%Q���x1!v�*IQh˴����W�@]] YEFg�[�8���DEԏ� ����|ǉu�x$�,�^��Q�<p��W|]�z�{��Z넪U���e�L��~�ci@����}���$:��-S�s�Bp��������9v>�n��R 3��i�����4���K�\��)�Ԧ*�쨥�p s����JD���A]��5E4m�J�R�(��_iykt�w���z�����]�=�߮���N���ȉ\N�J��[�۵�E�x9v|>��^|����GŇ��V	�}:�BQU�~�x�{w��f�ӛ��u=�ُ(�t�>ڊa������r�aL�"F=�}�.	1X�uo*��",��U�Tyʳ�TWLR�6�b'��h���\���I�Ƀp��Zv&C���<����)3�R^t��w�x=���Ǐ�2p�>u�|�(ׂ���NB�X�.�a�.p���Bl�%�k;v��&�$Ax�-�ǎF��(F������8���g����:@�Pl��ò�L����g�s��~��,���I�����+��?ρ����̴#��2��N<����Ҡ�_y7�O>�Z��ɰց�$�c�%
�)S��&w���y<�T�0zر����t�oh�;��	A��v��V(x��9�)��^S?��Pue`5c�	tR���'�>|����#n�����5�E����`l(��>f1k�2ϟXc���B1k�+!J#��V���X����-�;k�f� vMN���V���ǎg�@���1�V�C�qA;cP� ��� �(dh{8?��~�z/�.��,��J���ﴌQ��<����h�C��͵|otܖ��~�_h�!{�M�qŁ�N�_� ��S�Q�ݎ#h`�n�75�ZM-(+��}�S�rY֔�6�b��n�o������x�מ�)B�"1M�౅��������dm(�taM�U��Zĸ��C�X�o�6��g�I�?�ob/ v�B���iy u�w���:�
&{^���czw��,jsXڼ��t��!����&�gGg!�?����޺�)��}P��CO2�&+w?�5�,�������Z�2�=	��f�3�#M##%~�E$>Qq��Z�f?N"8O�<��C���r�E?I�ґ�?n��Ý1�x���1:���q�,{-Z�{c�V�:Mծd^"����D�� }"�Q�� A����I�GF��[�'�;{�gNa�R]MLv�»2��S�&ܬR��9���[�?�7oLt��z�	"��G),�����!Y$���P��͡��iƁ������d@�LYl�jy�8�2�hn�I��T�sL�ߦ���� "\JE�Խ�l�9:��-,�Ɓu�8��;��O������"�G)��t�˟0�RZ0&�?)�{�&yq�Ұ.�+k����0�#o-�
����U�[W!�ӿ�Q	Z	(���%��F�3�%����ն�=Z�B���Z���S)|�U,�[���l���0��t��圞��u�X�M��FϹ�[9�������v�
��7�bX�7��#�2�)D������f�4Y���#�o��{2,�H'i� '1�:0�;e*�&��a�5tPŲ�L{dpG"���ݍ�'��c�3��gӱ���MYYވ@4�W^m��� ����V�ȍnP!^vh���Y����@���֦2f��@b�q2�.�m��:�/���[��$$Qy�^qU�h;AoW͌Cae��y�BIM�#c������4ng�� \��KS¯�ӻ�������J0_��wA`�tX	��o�b��K@РE���}�~��zF-�Lp�2}����`ȼ�����[�K�?�S	4�ߺ# ���\��#����!�����go3���M�7���>��_N��Y*;��BE����g�#�Iܸ۸W��|C�������o��{���k���ve��F����;�o}:ǒ��j��|�@T/�Ż���	����>�B2��F)ؠ.{Z�2&�_D����Eu)���a"v��@'�����ɾ6�I���ܷ��!i�K	�F��/��:,	��ʫQ����/�"1���n"bk�� ��H<mD���y��+w�K�7��_�� Vz��[o��b0�&���#Vq��Uy���k��3��I0V�G��[p�kOZ�=���QE�wBr2]2�.�m���1�3��b�N:UkK̕�b���<�q2(q߯���pu���O*mhГ
^�"�-��P���M�� S�G�_����l�y%�>ϻ�-����x�JW'��J�.��&5�����(�dA��T��(|��_Y�A��";��b�>���NxY<�r���#՛����V�Trؑ�Q�����;n#Q���ٷ�R��/x�I3)�[��[�2�Who�:&��r��&"ut�Y8��5�KZ��ٲ()��0Y��h�碬&�,@� ��p��=�k�.C1��f�����Վ�
k\n6�B���J��/�0Q�#@�seb�D��Ȯn�㄀�\�{A�Ƒ t��b� 8~r5���;ȰR�S��V�m,xww�٩g_f����T,�y��7b6�n�A�q�:u�8ՙp�����
9o�I��$�#'' �q��=ܑ���`�bW�2 4�'ę���J��U�剚L�˫`���K�6�������C��]=6�o�l@�e�U�NM��� �,ߖ��������]�� tYRޔ9����;�����ry�J+�Rǧ��7�Y���ѹ���h����R5���"oޖ��Z4������v���K��@1��ېx�:�C�K��Aݞ�Em��D�.W�I��E��3�[��<u��ޕ���F������g/�t�1�t����.���g �"}V5�`3?'Y-��Q��*�ڢ7ls�4���p���j�����(S���U%�4�V�����������j?Be�`��k�G��^	��jCzh
joX̄�]<�.�M��+��2���);Ⳅ_X�Iٴ�f��J����%w3�1�7��냇�%�ܭ>Eq�okT�2�^�hCj��Qk���n�U�b�Q�#���{�4j�	�^@d���NR��K����y�������D6z><nhl���f�Z��9�_H�f[f�H�fHG�pAW�� *f��[�T������P����f�v��h�H"W蕉d&�|�|�E�_��d�
���[�.MMK��l���Rs�Z�k��dJ۲֗���.����\�j�*d�&�M>j�ܪes�l��A_AWE������~_��6�
����!�l��NjB������"��B� ���5K|$��[�1d��E��٨�A�dۓ�&�$8�
�q�$���s^��)2ѷi^-Dw�����&�zd�8re��a�L=<�g쎯��`9���	�Y�bo��i���">����dc�r 2���\@Y�cy��"�ү�G��_&��<,�!.��Y�s��r��6��4w�u{ 5RY&�TR:u�rM�M�h�.o���}�TrC�|ihjL	�&��邊�5��������5�Fs�Re�oױ����T��1�QL��<#4�rǓ���p�cJr�������;ѣND���K
��e5v��.�Wճ�Q:����*�gߟ��Q�~���w�3���u��}`��'lo�O���S$�&q�koqmEV�KX3H�2��Pa�3BۗA`��2g��4ٹ	ɈV��H�0$c:���C�P!nw��#��5bJO>�$�.�#��`�W7&�����3���4��n�x��6&W�F���0X�������Z������Y��Fo����W��7ہ��-R�;�P����1�?$rb��ĬM6|�l�H�/�\YT�(�q�3鐨h:z��N��|��˘�Z������[����3�U��#����K�'dS�`[@�[aU��8fuV}�8���+�d)wjm�+��� G���Œ�������Di�wB���D�t�iJ����Z�=�1�]:5��QgJ~R���+�l��^ �M�1����`!x�S��Zi���i��r�1�vЌ�Z��,��� �w8aL\��z}�a=���2��%/c�{п��w/�fãj7�1��c�<�q�!�~V�sF[��83=����'���-��ͱЧuF:��`µ*�C��n�|ZX\*nv:EJ�a�����r.�W�������:�
*]b��a;j���6�[������@C$�ˌ��bg�F۶���i��F1�"�5���.�P_�"ƞ��k5��(I��������S�/|<�b���Յ`�x�U�_G��UZ4؏�.|G��̔��L�R�dک��6m�������d5��q)*`d1��o-j��
V��}����F�g�^R �iM!~`�s3������z.V�!��U�Z�*A�~�`8�����ib��P�[��?U�2S��#u�,=��6���BǶ천��x[e�G��J�3�Y?^˪��m�]O`��e�8v���6����G,z�wΓT�kT*]hrfn��̑�ڡ�y�K���B�*q��t8�&�ӥ��F]a�~�BA�.4{�mċ�<�����}�sHr�X�OK$�\��y �*�~ύ�=���5����(��ZgA�� ��z����ۦ6@Ӥ6���^͠�b�"��#�I���� G�COv�ۗ�&C��^m�=p1�U� ��@na�a�/�ZL��t�����PG+������.����S�0�zU��:��v`錤M�h��CC�,���}\�*H�&�� ���+q�7�t��� 4d�$>=��jm~��4����g%���F��U`a_��χ*�`{��ϊ�!1ql�d �Ӿ�I�NC�J\=q�BTս-IDS�[���G�#j~���,����=<��ޱ�xX�����7n	��D����V-� q�շ��K�7�������4^�J淏(�D�B����y��ر�h[�(�*�t�u��]�p���*b�Q0|%=�%�Ǹ(�4����!�9)I�\[g�.��k;uQ[D6IB� _�o�G?8��3H�����iY/)6�W>�h��us��Q�4�(M+�H�Y�iKi��Ek(�o�hKD��S�nh�<:;����[ �I�D|�>��,56��3%v���k+�6�4>fmn�'�#
=� ^�����{F]�m?؀��ٲue6�H)e��.��d��A9��3��r�f(�vy���ooIR��!Uv��ћ��
c���D�����#P�="�l3���E �
Y�����fm<hm�n��է�������v�0��uh�r{�M�@WB�x����gl����YD[?�_Xl*���ł=��ˣOc��̥[k-����i
����X�ȟ*M��\ǩ�(��%q��8S�K;�v���	c��Rvn%P㪓�d�i'J��Kl���o�������E��6��7�a�n��	��h��vr��to4 ���w�U!]��Ŭ��M^����T7�g���k��x�l�c�1��Ϡ@�7;+��9^���Ѣd�X۷x�̨ɲ�/g8'+SQ ��n����p?
���ժ�Gr��ϖ"6��p$�7��b0��ͅ�����n�%S��L����垐�ۃX:[y��I�g���3+8�s� 2�3E�.�L�99z�H�^�;��^��ԧi�b�<������EszCr��9z�gc�����b�dJ��{Q¤�n����=bK�H��XUږEk q�qۀZ�뼃F¤�����x���+׾�RE���\�ky�**rL�F{�he#X����|�c�����	 ^3���d�Y	���(;����2(#ǯ�V��qh/�H�Y��n��ܲ#)�[���ߺ��+�)XpZ�0��qs^(��bb����`��u�phsR�����D��9��������(;Ⱥ��n �f}�7�o���i)���bt>�^��.�	H���ڼV��j�*�8z'aj\����`Z����0#�5'�5��7;��=햗s9Q�oc#��t^n�����"�1S P3�
a��4�o�;T�1i�}8���z�v�O�A�µ�A�� B��T��Pͯ��Gd�73�[oc�l�L���S�'c���Wnh?�:Wց�J�!Lr�6@�}�y���0=ҫ_kL�y�x:t�5��iնLf�nqf�I�����p�߬W{���z������c��	=�[}��5� r���DL�Q[�����=��}��n�4�6�cyiJ�U��u�O�0%�f?=�PQn,�/o�m+�%�,��,uuiZ� �q�)c�ƻE��>��4-22
�<5n$`C�%%R��H��,Nx�[v}F>#��akF����{�Oh������ȝ	���f��>f&JZ��Vr?�H��rE�m�t�r�;" �_��_m��q���C�*S��1���%ٓ��O<>���~���8؟��m��l�IR��r�V�<��Á-��������P.�����?�t7Fl��$�I���Ŷ����bޖ����S�%,�#���:�&<c�G��m7(D;��a�q=�T=�p1���<|J�*� b7��e���޸�͒s��	5�GU]E(K�BP�P�|4�{sU���&>��+�A����<px���(]�(G��iB�Y^ku س6��'��,�'? Nt�^�L����+2gMD �ޭ���hE��5P��6	��C;��{��5�m�UiAT��G}��s�Y�7������:X]���?��NIjcri[�\Y�+&���u�WY��ŤK{��_�8I����wZ�?Q�Hf@����AW(pٯD��r��P�+^�����v�l;'ՀP��kx��f@d�R���r���8�i��8��o��V���c�����z	�Y_�<}�<Oݩ���?��YyT���ŒL�|�Mݞ'����Q����������9>�/rӐz�Q�D	�ތ�;]��w� )-1mp���	�773�:�s��EvG��|=j<W��􃎥(�Ʃ���<�b2S{�!0�𐦉6�M��,skX���gz���u+ƒ�js�!/?⃺��],N�}hu�x!���ˏ�ۆD����C�����-�{��섨э[l�e��W����X��κ���쫲��|�����&|`��c�"([�����		L܀Tv�-�Y�A�ps3�:z���ըE����'޺�FEDx�����;A^Cf��b�KFg��|�`�d��7��à��6��	𙟤vr�*�u�` ����\#l�s��T�S@�|9�<��Y�`�����l��!b ���%���NBÁ)`p�E�[��?��ϥ�C���-h:�@�0ާ��5��S��6F�~m|t�c�� +���U�$�_�e��T�` ��Q�a��(]p#.X(�{stP��\)L�Φh(e;Z=���M�˦�4�SP�B�/�tۖw�S������n�}3��l����3$��q�Ԇ �N9x�R�$"Z��)4�Ǻg��^����Ð�Բ��4���?t�rxo�3͐]�T�ߟ6��s8��Tԩm~�!��}���o<�\��<��&�R1|e��y䇰��<T�t��\�:j�Y/:�8n���گd �y��I�(�`l-���R�Bޒ�3�מ��2�`�2��đBEYG�B'�DgfK{�r��s��p���T"į�甎?�R%!��� |0�R7��;}."�]���$�����|�Z�8^^?o�Ȋo����I�G����]��
X&� 9�2_�?�~E�;&�$�5�i�b>�-�B��_��l���չM	a��o��!K�.���]���,wc�9v+*��؏g�=)�+��0I6�S���}<#�'�g1�����1x��k�Z� J�!t��xo[������^n�����7-Wf2��� �_��;�i���/����sG�}�X��፹��U|�������ai����'��M'QJ�i0#�������h+�+�<�y�:�����f=�9)$q��	q7�ʤ���}l�����<�^AĊ~��1�`j��:�szXD�$���y�3q8S3����n��#rU���u�Z_��EQ�í����؃bc���ڲ�֙��".ɭ���� ���u�5y)�%��a���Q;MW�{�e�p�ғ~����.&��Y��<�6�"e��ʟ��N�̷��Cfa0.m'���#q?wuf٤vp
D�B�b�'K`
/�π9�I��O�8�)KX�DqU�:/������Hs�pu ��_��P�v/�n0hp@�C�5]߅����z���D���FI��HĆ&��'x�K�ѱZ��W_�����>�������M���,��;L1uÊ84�,��PC2�{��w���MFo�Nw�$_����}��xD>�Y��+�'Y0�"���(�D�~�����-X��Z[������S�mq|Ť z�A1QX��vK��@SOC���dqi�#}�_��6�����Jm���e��r?E�g\!K�`Lў��>�O�̢��E��ֈ�t1<1G�ޗ!��2�t��z�@Te�L���#�ZX�TY���������T�|	�p
� E�J^�l��)�dx`�X�w h{��x�ݜ��F����Y���O�$.�C��4Ӏ���-8~���n��qP��<�;���7�g��Z���֪�Wy>h���pZR(��ja+G�OK�#r�_]�0��;S4���	)!,��m$'d�S�I���D�"��4%6��-(K����4x�D3�ZA�*��a�`��%�J�r���e �p�Hh J����_����{ܲ}>��̷�QP�d�������چ�����Y�_Вt};���)it�I�T�*p�(mcv���4�]��`�q��ߏ���k�]�͏��t�rL���qRz� �[i~Z �'�b&���:p��r��Jۂ�s��;o��h35U�����y[��3�~E������!f,e:c��U��m+�[��Sa-��+��^��9�QjP���Rp��G���`�o�S�BW��RcqK�2c>2�_,V�6�E�o�5��ʓ��V9�<�j��zoV�׸A����ʱ�IT�y;��S�߅�#z�ark�w	���Q��+At��O�y �m�W����y���y��Q�[Y��;(t�Юs]T�Y!
�u��X�a}#n���"�w�j�Ʒ�M06f3ՌF��D�C0�Z&�ꖼ	A麕q��� ��"�?a]/:k6���B�1	0׎Z%�^�kb(�a2Ó�t6c{�D�����5�	��γn����%����T�s���Z�L{��A/ځ�1@┌N�J��!���"����0��$�n|b��5�#N<�����y���E�Lü,��`a��-o�<���2�.)�z5g����3�H�? F4W��!ހ�M�����g\g�F4:cI�g��~�$���/��P&���F�5uT�2�"�J�6�|�����o�ڟMq��9�������k����mZܝ>�h��˶2�Pt<�O|��yNҟ�ۃi{��$��k�׳Үi��<;�"�*�sL���=��cU��{6�9��H�ۯZ� �k-��yd�5����C�<s����:�"��]���G��/�ԢL��G �My=�����@qm�8�=�:����f���k{ �2��?B�����?��z�r�}��i�2POf�Xq��o��U$�3N	NwB���'=��G��"(g���B{@ѐ�/# �J\����*]q�_�f�1qsRv�����~���q�*��������Z*6�T���@+��⢽5[3v�S�Y%���/
��ׅKq]�>D��[B���+�=�{��\�w:�nн#ɒ��ݶ��,:
wlV@?��,L�
��:l�sT�)�����ٻ*V^ ��@��Ȟ'u�sd8�D+�jW9����!��Э���#��� ��P��hq�@�X[n�S�1�g��0��UBM]��@ӓ
�x}�o�[i��S�F���#j��@s�%/�*?t��WkC�Ҭ��٪s�M�>�(\4Uӣ��"��w�W	�j�7�W���}k.D��	�,r%P����hUD�=؉��^�����p�����kO%x����\������6�n��2 ;�N���xzX',������,�!\�e�B�T]$FiS��=�����n;�狥yxy�;`����g:/���x�$��qX���V����Kq���[�c�
Fb��&rW�MR/wA)xK�(LT���*�np�Q=}2L
X���Ӎ���Z	�O���̙�@�����y��@��9� ���n�
0<��66X;�m����