��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1[@�"s`_�Z*���Un��]H}k��Oi�'$T��*�k��W�B�r|wUxED`�"��&�"7w	�Q.e(�el�ӿ�ú"��VȠ��\�&q��)�$�>F�����t�+zH�E�(�H���O��C}�y���l�{�M~l��	�=�|�iֲ��,���� ��k���A����wɦ������7���or �ܗ��1�BÓ��=G�y՝�J�kDXr��QB��?50��b� S�ʙ�I|�&���%�M��x)�����\ �J��|E����U��Ys���`�b�@^�k`�K�#��5�M����A"*0%���7�L��t�M��DĪ�D��OYw]�����!䚖~t��@�f��c��b��0̸52���6?�ˑ�²
�gH�ϩ�zQ����ո���5��}h[���:2���H�Kġc���'7� �+_ݽ������T`¶��Mt"f���8���;�Wko0D�с!^I9ƶ_t]��*7W�I<���!�W�ܷ[�U��L�>}�:�M�O�J��2/���aO���S��f����} U��GS�P�0):��>?H��r�G-�0�����U`l����υ���]0������0u*'�\O�<և��I���a,�8��r�ǥ`�}�SN�f��+�]Y��m���`&t�W��5y�bx�u�f��(��	�'ոr|O��-UㇶR��0�4o�T�߭J�t@f�l�!�85��v�i0h�J�M=�qbr��Ga��F�S��v^��&�/5�n�_M��9� 5v����,ZK�c$��x���
��Y�����M
���|�@�v`��5˷Ƭ��a#���R˴�@��Q{)d�n��T��3����"=y3��%�\��I�Y�=���g�"�l�t�2�]��k�S�u�-4`'V�t]���=Y��+Nǰ��/��Rn  c�}\M� �*9;��Q����RAR΄af��Xe�K��ڼ�����ǂ��E��Xel�S�y��w��}������2 �A:�U�oY�}Ȏ��w�.�X51��n�`��"%��?(_3�d\w�l����}K �Lf�6=\k�
,*��^�4zÝ�N9��M�-�)�K��P����VHY�Y��)G�m�5z"�'�Q�dt��	����z�@�l�KP���~��=ic��0�Z��`�����&IYj�uƞ�MN�E���C�y�Ш�JA�nH��f�hXT>�	��X3bҿmT���is��鿯9D�h.yO!�t���弃����bJ%�
����w�t��)���R���F�"]������
�yI*]�95Ļ����*ͿCiö;��{��o�=D5/�/���*��,�Y��
�5�ZP&�Z2r���c�k	'�X�O�␛��)v��t��Gu�Ns�`��q�E�>Cd�P���&�F���,��V�R�kǋ_g%@��g{P�81���$�bh���~uh������8X��&� �Ή�����ZKz8ۑ_�p���|1�	��_=7 ���X /^(������*(�z`�5�	�?����$i�Q50���H�v��u,�_80=pu����}BE�W�a�+�)O�R����i���F��~���b�B�����8 ,�C���n{��̧��&!-{US��9Ԟ��,w)\��K�f%k*��Q�U(�j��e���U�?]N1Ue�\0����=����P���V<u�0����o��t�;���ª߉T�xs�]��ZX؜����	vO���՟� r���9XF�{����X>����WH�#��K��������@���L�A�_�(�,]���p�',�W���Zt1��ic<���."�U�N�o;)HG�q/����'X�9&y`+��0�Ϋ`oh�h'RӝPz�s�����y�T��4�)Tx��C�Mݜ�I�O�W�-b�2���놓�m:=&j<U->�䙣�K;���1MG`ah^���l4��C!��)C^__d}���?��*1g
�z�5��L�+3�g�`�%�$k?
z)��s�� �1�g7�&����NRߩU0�4�f�,�ϕ� �lL}�DL@b v	4Y�3
�_��좐��Q����u��P��K
<jN�;�z���q��JlZD@�~D_��ԍo�"Z�j��e�I�Aʮyy��5b�Fw�+Ψ���~d"��i���w�?�Q�sP�)�1-��X���޸.��q���LI�`n]�W��`�b�9���;�&U�f��P8��H�%�uM���Tt�����>�HT:<
�Qgқ�V�\��BK��G���d��!�"�DK_T�r�Bar�灸R�B`N��ʊ ~�!�L�)�ϿPuR�luۍ��-����1X��i���~&���a���x_`A�s��tʛ��-���*d��O�����G]�$����l,�D�T�4�n��7a�wQ��|� ���<���*;S5�	fI*6��傿�k���-v�7p^�}�:Bj��[X���4���a���sQ�q���5o��/[?y^�ύ�٥��V=�ڜA�gCXTt��	�H��1'GoW��c���[�v�l���cg�BW��'8�.R�����zZ���`4�K����o�=��L@ٹ�N��RQ��`�]�q�N���X8S:�&C<�Ö����	%��<����3�Z���tV5���ƄG���趘e���\x������Q�]� �����a$����Wsr�
am
| �D�B���3�E�q ���r^U|�'�I�0%�z7����*��#����!�h1�m!?1,&��T7A��&��H��R�
d�9���2�D_!Q��1�Dx5��0��q�Jd���I�!�Ly�?TIԡ��9������b��@V �#�#x4���u.|^���\e�$��9��~��P�;��������|�ĿAj��۵��s��x��DK�|�&�PB�:�}C�Q��XY��H_1#[H��'PH��YG߸ܫ�Z�����R_�)�"ܨ���د��>|�՟�)%(�q��+q��v�����#|���w�Z-�=�=��&TK_yAp4F��w�ֽ>��ХY��(�eͪhߑH���VL*��?DLԄv�w�ipl�O���!ؕ�c��v�9�����;2�^��8�?�PMT5�����7��V�����,v�[�t�����Vdb�K9���r�g��oqE�~�Zv�/�mʛq�E����J��ÿ�1�Е?*A�	]�T�
�F��Fv ��2`���Gf�I�P��!����5���v�������)��◁h?�	�������6*��EbNJ۩̦�ϒ5�he	��E|�:~l�ȋ1c�o*�����2B�'�F�ڃN�����2[P�v����	O�����%�4�� V�J[>t5N���*9a���]���,dw����p_	�) ���3:���V;�n�+��Ɲ�N4�ޢ4!�]�-�U�VE��۫r#���n.CԈ#����`�|�y�J	jF�eer�B�9mgV�,ʼ��P�̸�SS���ҨR�U5吶�l���� Y�v2�M�`�S��h�N��8d�ςLͨ�˧�kTƗ(���� hV^���'�,#k~IR�����>U��Z_�~���<S�H��YE�U��"�S��T6��#٦�+�������P�u��ڟ���?|�bx۟�3��t��/���Rn�)��g^�,��2t��f��J�ߝ{0��I���9�q65��G�:�{��u<i[��`
7p�>f���d�'�kRs76i��|Ο�����4ٺ�ߢT4������:���&��#$5�z�83�_��oҸ�T�R���`����$��G�����аDT��{��y��%�X��=���'"[���������@�H�S�^]*z���ߎ�g�J(�p4;��tT<|�����A�%��(\|ө�RRҀ��L"
j�0/��6.p
�.sᑸ� �t�ѷ�a�ظ���'�I�$�3l������	�+4������p�l�Ai�T[�6��a��Ǵв`V�$��]y�!x/G����u��}���g7���CSV;��F���&֑�m��#3F!aEk|+�)��4v�I��4LPJ����Êg9�>S�ڃ���݀��Z%���f0͘4S(���V�Ո�2!��i7��C��!C�D��`^��^��Q 9H^�ܚZ �U��KPrlIOVJ��;Si
���~�r!������|�X%�G;����$)Ju��8,�W���] %�s�p/�Y�WR�q�,����_��A&%.�|[��L�Y�0Kˢ£�5���J}@~Ẵ+/A�Ed[ً�CF'��5	�V���b	Vi�Ãz%� <\��?���Y,O������ʛ"��!cQ��T)�H�ގ��9v�Km��d)^o۝�����51��_51��3*����ZY�e'-�֩(}��P��!([�fh��=l��1�D����C����i����ՙ�ϼ��������+�[�dJ�w�k(4�����2�rST��-��y����aCF���7��]Md�D��0%	i�v�i�Rc��W.%��m1�G��.�:n�e��~U��%//��R�k�Yߠ��^Q9�*�g8��4Op��D����f�EL�Sސ�2�"��w{Q�`�5yC4��;P���N�5�.Ӂ�#BaYc�d��uqIK�V�N!����yF��Tȝ�B��irddT%䱑�a�A��ŁƩ���r^�Z�{>��5m�﫵o�.�A�x��%��Gv�"���S����1ٞ3bF[�+*���#e�;g4ռߝ�Z�M���گ�6'�x��>�w��yc��S�M/E�@-���d�S�2��NT�z����WuN�M����[dy&Ff�%��r��;��"��F�Y9�^�e�B�=�=���ƙ�
��VFD���^7/=ST��@�b!a1B���2�&C�p6���y���{N�X�v(���]����@>�HN����[?Ep�� ��Ʉ��凂�%&C��]�|>وJ &>��.:d�6��A�k�k�I�6�/������qrƴu�ͫp�����T˰��`���Y�XR��bt-�k����R��(�}{Tuα�z�;NQ�n>V����*�6ٙ�_�I-nD�l����W��(�/�ן�3��G�e�5���5w���>Cx>�>T{=�/ƭ���ʶ�0�w|_Xg��yTP�۳ټ����u������U�8��e�G6:�&��b�q�-_���w�g�|=O�;�N_�c�2/�̿����ؐ�=��3[X`�xȶ�L{����'T,M���q]7[���Lw�%����5���П]k3�tp���n\U�KD?q&�p��*T�*`����b��;k�IE��u���lpх�Ծ���I�J� Z��#1<-b���l`���(P�Z���Kz�m`�>�!��Ե��h�t��[&�Wzw�طb�g*������
�Np=Q��9��lzY
���\��>0m��Cٚ����6�\���R�9�X��Zܺ��+su�7]�xKI�L�ɲ�5�����)G��'��r��d/ŉ�
 �-��(BL�'��yx�������lu�5��]����ͦV�@�>���m�Bq7�Y_B�us�xyg(P�i�1"W���ԣ�V����ܷ�U�h3�9.H�v-�Q�X�ֿ0�'i�ngDzt1}��R�H��ՎQd���dU��'�ҷ|�=����mġ�)H�xc	v%�O�Ր�.L#Z�Q�0
|o�;/��:U�su��!E���X�}q����,�M-I@ì��#���*���k�O���umk����.1��,0ű֜/$G��h��;����J��2�V�S;-�Y��r���)�U_jfuk?�j����;��c(��;HV���Yl4��T*V�'��?���s����5F�݇I���=r���\��r���i�oKog#0�<�[/W��M�nGΌ�Z	w�<ǬԚ�к������Z71܌�P����"Ĭ1e��xSЄ�uM�/���/�j��2��/�N�'�-�̜��L��M��2P5��H[;�+�wm�Gْfy=����h���_`u'��7҄�~�Q0���~��yB���M������ǟ�
�J��J_��D忬�M���_�6�w��-9+�Ő��-UT������f�
X�ު�|0eyu64Ʈ`��}d{\hn'��ĮV�Y��u��	�u����`I�hN�`~�Ԧ23^�ڧ�ݼz�vg�7�x�<B��eseV
�
d��hhUvK�(���FH�Lm�c>�6	䌻���{����W��s���D�pd��4�[ �}�j������2�
�����c��J-T83R��Y�,�&/�i�.��@��O�T��	��u���>
Ůf��՛��"M��~������a�p4���4���f;���r�A�bK���t��L:�����{`"QVH�l��ϩ��{UVne��B�.{�*�񿤷����>�b�:���lƜO�5��Z2���\�8Tzu�]Qͯa�Vr�a�p�<��i�X��ftUh\�8j�CD6m�:�Ψ ��6x;�@�5��7�N�T4�J�RD���'p[�.BA\̛��\���.{�w y�u����#Lة�E�H�"*}&qWS�6�^g�e���k-�r8�j"��OZ7�k~�ֆ�ȥ3�QƷ
�\qq��,�lk��o�@P� �_���O7AT�B��\�U���������z���'���ǅ�_��7vm~~�z�u�YLLA��W=^I�/��ؗ.`���$�2��#	7�Y�U����=5�c�gTYlF�u@�5��p��K�8Vt�ߝ	��������n�	�uā��U �J\8���gu%wC�&�K�q�@]Ǥ
[�?	�&����h�� 0��.�&�����f)�Y�M�m��KS3�������hc�J���u�T�ŋ%�@�s����B�ݞ&�
�6������J��6d�	�'�l&���"�_ZcF�U�٧��1M��o�8�LNf�c{wH�#
�jrj iq�0s��5���)�'�����J@�����)��7�p��~�2��KY��}�'nA��DAd[3+49�1���Ƃh�
��Z_��h+�Π��,�rv[�ſBGߵ��=��$r��:� Ԕ�O��(��ڒ�k�S�l������fX�f��Y!UQƌ[<P���ѫ���h����>��X70�ZzJt�c ���|���\�_5��W��}�K�����׿�y���c!����)-��g�rp	�z�� n�!�~���G'�g��.ʹ}���V�e���$wqD4A����$��Xd���G3�D�Ő�F��G"�@*iXzW`��j�V�!�7�����a!��S��r��VTD�.��*SZ��!����4E�=8܃`Lʼ���H�uUtU���@�"әF�iT:O�iy��c^\a�&���!ah �䱞*]�<�!X�R�0q�pBd`��w�$�P�rd��������)��K�`=���Q9 ��l,!�}�J�]�p���ʬ6u�Ol��o�N���'蓿�͠���k,�=���d)�T���9�p��uY�R,�c��M�����7��)xF/���H��⠁�jgAϞ�#��R�)�b=��6sS��&��.i���Ǻ$E�C�`

 x2�z)���7�-䝗k5
N�T���-	T3Ʌd!s�ln��e.b��Aw���������K!��� �fhŕ�����*V��N���W��5��U��-�</r�o�$���aq��I�\m%�I)<b���қ��2D��Di��L"��b�[��k|:��q�Ձ����Q�4�X�^��lY)���kz0&�`���|]�������}�;��� ��4lJ���ɶ�i� PK-�v�z|n��.���0����c��w��@�?�ybh�����jX�(!�����Ю�y�yo�M�_��һ�U�m;������3I������MI��9�6��3B���nY_wD�z^*�]C�/�;b!����SX˟��tsb�B���#��:��h���,?eȃ	l9�Y�g���_�!�;�=�[��]D�f�����~�}	�@���Q���\[�M��ԙ�n�WP5J�P��ݳ�5� .9����.�˄�&�q��N|	Ol�����`w�Rt� �K�C@�.%�zK��Ŋ� r�(��>ձz&�7���fY�v�뜦6���æ�`�����+����U�1d��{b��`���'�D�`�i����`1�fN#���{7���c�m�h��Γ&W����K��7������Km�:U��4&X�BDL�P�ϩ�T�cJ�k-=��ODW��f����Nh�`{��z��I�]Yۄ��w�w�eD��xF�j��|B�Vu�5lM�/|�v����I�2�6�ʯe(��6�#~�h w�	ڪÛ�2
�5r��
H��=�(9�?@vWlt/|����������u�`�v-'�A�Q�%�i;�� ]�֢\��Ƽ_E{"P$�l�̦�*,;����T"gwA�Y{Ŕ����Ks�*C�0UK�?]�
^�qy��Έj�gW��r����ܣ
�Jټ	�A`�E�K?�~z��!4���^�%��U�3�:���Ls�vC0tZp5Y�,�s9@d�~ݍl�e�����hW����׶'1�P����5�~R�i��	��v'�Sx�CW�jx���.?Lؙ,<͵ן[�=��{�� ����`�����**�S�+dw���Uͅ�x*q^s:1���(��Ӎ:ܭ^���YK9�R@�h��Ϙ�\����;�l��Y1��Y��6�#�I�Z��V�����ܨ�?>����,d�$)^32���w� N��鐋�~�_{�d�ꉻ��  �|$���I�[���x�_��܍��1E[A�+]��+�'%��\w�V.ߥ�r��H�x�.P���v�م���i�[K
�� a�2��6Ua���m&j�%a��O%�1+���XF㎋���\|�׎x�px�T��
 �X�c	�~��1����jN�:P�a�ƪz�����)ܵ�,1yQ�SmK�T;��y]�T��p�#�6���W @�w�ѥZv����4�����qWM�B�?���Y��g�߈eŧ<�#�ɳ��<�}��3���Ԓ�4'�(�XA�����T�o?�d�l���:���
香I���r>�JV�JQ�_,z@�V���mv���F��8MR��7�ڌ�ݧ����U,H�b�b;m5ҏ�02�t,����j>�����p�)/,�]�m�C��*	 �ED�S�?P�#;ac'�����c�O�Ƅk*����/i�������4W��UBf�%�����a�̰��^aţ��o/³�w�QX�{d~�|�@��' �B|���m��� Ӭ�	�G�ި8T��O��ȼx���'�*z�A�ҦK�es:B��4"�R��8�ʽ&г�e���W=!<?�
f��6���w"f)fNuB,��ѝ[�����L��0igYZ�^O`?<[m:��sԳ�v��B�'gB��_�M����P�/��i_�x�����fC�~�%��3��j#���*����wf�Ѻ5��tU(e�s `�5\����r�t�!g=Ti���>XQ�t`��jH>R�A.Z�[EA+Js�� F}b �,��L���~��/!1	�H��{3�uk���9�X�f�T��x��D���q�F91�g6��z�q�?mL�W� t�C�a�vK$'���7����v$�Ylp4{�a�*)����09P8�9~�o�We����px4e��	�d�w�|h�W.G8��N� wCj��bu�����N�>ꎟw��]J����]�Rv���H�l�T�C��nE.q���J�����ޟ_�0҂��@[5ҭ}��k�j�nN�'|T��HQ%I����b�]k�P;����2Os�'�#+]y�7� HƇ�ژ�<��rC�~0�!n,Ř�����S