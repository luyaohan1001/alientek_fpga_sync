��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ�;+G;�2��\���|�Z���hX iK3>�P`��&I40�-z(S���喔c�K�_�<�=�����
a��B ���������w~��t��3�I��b�Y�,
2s���b4Q�0�?ۯSD�>����ux���.HG!5���p�N�r�.v���o��;���98px���"������+���f~����"]4��x	b���$����R��s^��4qsi����<K(ǯ��0�^������s`/qO�ِAQ���fz����
�Gڷ�SA{��d ��d!#W��6d�v��x߀^�pE�XdTZ��{�΢����#�Ꜥqm��є�!r�z*�<����(��� ��Q�:of@��iW����ב���劢�%\Ŋx5��K����״����)���h��lo?�*<���ɋ�G��<J��N���Q��@��:�$�G���ԟ��9��2��NA\Țn`���עx��X�<�V�Ȧ�F�Z^ó98#���� ��a�B��c�S׸e��n��e�DY)w�ƞ}&J^9&S,tս�6rJ]9��oHZ���5x�,	nH_Q0ǎ����R�=*b*X�C�]3>�A;-lʈ��ˣ��h�H('Fr�{0�0�c�)�Z�#s�h���
l|�4�$���&�����s�D5�ڜq98q����1�FA��ŅY�dӁ%�z���x����)g;�{WF��Ӱa��O�$�������^b����EU|6<�ј@ڢA	��KQCT7��ݺ؃Y�[�&�>��}�$��kf�#OE|��	����p"�$tՑ?�k��e��~�.���&䔰�^�lFYAɟ��.��]���s)�����C���WE��aR�yj]�	��/It��]Y���!���w�0�ࠩ��ț�)�l�5��7�BLhIڀ��O;le�_*�S1�&�5�c��J�T�恜����\ܥ��K�(���Q�뭄%L�+]
p��Ft�5LTk��`��xv���3�י�\��P�zƖ�^�O��[��x����T�}�( m�	�7O�t���}��1HBа�8��Ef��>+�f8{{�C���q<��Ut�����&�4��i%������,����ݝo��������:0Ь��jg>?U�bN�4x�pҭ\��}x��&��"��g�az�3Iy��Ԍ�E3c�o�rx B�q��A��A/އ��:`���Z|/-B��kJ���71Q�ڀ�ŭ��:,�b�E�Ͼ,�`)w~�D�D�%�g�$0�B4��" �2z"�PWjb hr���ItZ=���خ?lU��0d�Dl�/�S����6w��d�\А`��p��p�Of!/k�Y�I��%����P�A��\G��f
��4El/`1��6,+�%\T1��$qEIW�B�V_��R�:2��=�4H�*ş��� ��c{��w  �'�aG��=�9���nwp��f���'UwJ�G���;t�mѻ������o�Z*P���m�9*
#%z����K��%�#cWJy3f(�q¹9���I*�$�3';����a�!w�6d_r�7s�;I��IS�k4��5������ZZߜ���ԛ��Z��<#�����v�M|�]�3Q��G�v;ėʃ����eP���w�9x)���ˆ�c�a�3z�ұ6y�#�Z���]#�
�IJ�������sF��̬E�ɩ��-C��A&	��^��B($��%^�V����Y�ş���vxX	t �Gw�^$����s ��#����O>E��y=y��&H4��z�5)���$ϼ��@�R.i��v�\�-Աau_��7���]aX:���� WX����X�M�q<'�M�������z�4��^۽��檩Y��*V:&�sD E�KF��o�Q9��7fM�Mo�fB�ΰ6 �F"�eu]�_���H���.�t�3��0X��f\�.�.N�⬏���Uf��