��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL���m���C6%Z���%�t;E��QZ2 K����b��鼊z$?��ƛ���V�W���'�(�ilP���Iʹg�f�����u%@�3�Dfc�PDгR�7�8���E[,�:���*"O�L�/Jx<]-�Ɍ�����S6�U�%�FdLxN��F�/t(w,�Ú�T�n�����'Õ$�%�4W���Xy0<#��'*�����V!n �[2:3aw"<rK�ko�f?���57o,��[M�=�F��Ӿ (�A�F�V
�ʖ~��K���a.��&��/�N�=P�"k$�j.=�
���-q���`�y�=3�$ՎR�9ʲ�϶�8�O����ayǶj���с#��n�����U]��t���*�C_=��Y��=��XP���l�����T�=�%�7'��]/'p3b��8�[���
�Z�e!�K;wR����=I�Y�i���^Չ�U�(/
�bx?�}��J�n���7JJZW���e1K����`��uwR�~:��;��,w���y��O6��og��w�mQYh���6��3d9����H8��]l=�a�$eJ���ȃAft=��Kr�+&b��ܬ:��|��VB��U��vz(������5�m�ݾ�Z�<�7co}��wm��{a�8�V�`	\D�'��G\m�r�[�pl�lo�f,t�̛������)V��ͼ��UM�=�a!J#��f��(**Ρ������+V|nC&�)>ti��(��L)�~'��4�T/q�b���Qk���|C?RNe��xL0�S+/S[��M�l�j:E���f^@|�2Aj���p�k�����T�����@��ZQ�ҳ�wў��n�8�~��q�J���E&tRi>�ld=�r�YCT�V�Bn7�^���"���|��� ����K=*����:�9'{�]xb��i@���1P>���D�)�}^�Y�<�(�0-̻������[w��/�~:���b��}���U	Z��D�Y�
�y�^B��VW�%L%�h���V�%	x���i��B�q��Z98�����x���mTĳ$�d��}�	cT�����G���ah�7}�����-=|�w��;��^�'���1g����%B��p��z��(W���X�x�Xӹ�=�"{��`�٢6��R�D�([�W$���p��Y]x�z��"�>v5�5G�9Vsq�֗��k�v����[~����@F���W�qxC{\�B�z�0���_����uE�DY�G�C��l<�!��%&����v��sj5M�$���/Q͐L�/(���m�T�;uAS&�{��ٸ��/�����m��9v�t�g}���:ОM�ڨ.vSKD��ˍ��P�y��YM�i�@8'�B>?���Id-�oe{�������]�Iu�r�3��;�nC/"�,
��tJ�`m�`��i��#�s|5������
aR�S��3��HIZ��~-u!�K���=c��\�f���_}��+��&��b�k��y������+U7D�䟸������d٧Ah��b�Q���#1V�q85���k�^�Uu��#����`�5���J�۽�?0"�jO^L�T�"m���"���릗� .��M�p@�-b}9��OwT���p�:2���'�70<7�ؽ�cHxm0ˁ��{n�����hu�B��ӏNY�m��Z0fʫ�������=���E�5�&>�
���P����p�w=�k��j�D�EpL
R�Up�����P$���*f����_�dD���`��LI�K��+c�F3�P!6����<Ȅ�s�.;����Z
��C�������;)#"$^,z;�e���-�սN��Zf!��[���j4R��4U�0wܓH$G�?x�A���EmK�:!$�|a�5��$(��#{���}�U�(B3LJ��>��3`�����uC�?X'�xq��
-��Ci�
T��*͹^1f��}@��r�a��;v 8+���3���fQ����L��µ�XAH�O�?�!��f0x�H��Q<��Q��l���6{K������2`��*���U{x7���:/�٩�!�w��X��C�� +Ɉ�eZ���D�@��䶛��FW��)F[�]m�>T��je���4�w:��]q��t��/���^ ��n�1���.���WF�Z�QQ�T���ߏ\���L@7�s=.�}j%�My��+B�|D�8rx���˰���sXT�drs��M��8�-<���XqO氯���d�~��3Ԏv��%ZI�=-�ڧ�+�14��Ì�,C�5�(�h�Å�����W�Z>���yަ�Qs�� ���)�#PV5�Fh1mF#9�\a3�;^�6��Puo�.H���R�Ֆ	p�ʰyO)��~��KM�]Z�Z �6�vB�1�/��Wcy�
6Y�����q
[���!��Fn�}�|�x��'p������L�2W�y\�(�e���&�Hjt����N
��Qx��<J��:>�+�U���n�R��@B��I�\���D�xT��ۈ�����>R^�R(�J��d�f��فoR�)ꤻ<�|[�M!D;�ܣM*Z��q��A��l��"��Œ�7s`�FBl�$�&2YD�0N-s���m�C6�}(��cL"P׈p�g��)>����Մk���R�	_��聾��;K�m���,�|��$J�y����e�(chǃZ9�O���R�l��s���ٛ���#{��p���ق�0��N2o�h�$��1SSN�4bӏ^O�_G�J�Q�FJ�B]����I�n^E���vT{+ٙ��`�Ϣz��f��__�$
cՊ���Y��7����(ٸ�i����� ���������K��n�J�Ğ��!����W�r|�R�!<��)���q�F��a�����T�!;��]�
m�2K��/p��U5���ٛ���JM;�}�^&I���'����#��K�4��|�4�=���?)r �j�^iS�+���r��\:@�<��������(T̃��S\j�����	���O�4��P��L�Ჸ�9X�=9 ���>4K{n������i*�B<��`�l�I�;$��3�kB�_���n����ZQȊ�A�I��>�Η���*'�q�vY��V�߻-o���)���Ex�A�ۍ ����@WL����}�
�8��~g����$�n�6����)[���ॢb��	 Xsn�POr��BF�Qm�o��� �L�W�[t�V�Ɨ:O(�"��s����9)1 �]ڹ�rq��
H���H�T�6��\\u�����(TLY�������vy
bw����%5����R�x3�N���