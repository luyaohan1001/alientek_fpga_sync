��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL���m���C6A5#v�<���B�kV4�74�ц��M��	�e��:e
�H9�GK�62���U��Y��s\���S�l�j�q�P�q���� |�M��[ġuߚЈ5�W�'����01ָ�7]�����˩�|}D*��7�-g�B\+�`������]7�繯�QpxT0�'���֓�G\!��d"�u��6��i�%�1tIv���q�6"ۅ26��9UgB~yB,9D<�o���O{Ć�?LG�p���k�|��,��*I�=� �ƈH�\�0-��j��$�p�	)^ \�}c:,|��{�%o�X!���"���?O.z'��N)�s)���ڕ�H8(1��2J��)��u0��n�v��"�������@�~�s��g�j�����^C���-X���:+���[�����U+�h�ꆳ̣s��B� �>��b6���咎s�3�y����I'r�#�z{��Zq�P�I�B����=I�<�#���=L�\PV`&�Z�uÒ�f��O�/��]�Ha[#�2��
�/�"���)��D�#�zL6w��N�k6��=�X�T#�j�H���`��J/�c5wF�oO{*�R�oG�`'�./�"�����jDm3�z_#���U?��Ne��f"|/�f��%l���-8#�p���)f��uBj͊X��86+����J;H��	/A�dҡO˺���7٢X1$SE4~�L��`���ث�	� WXq��j��0*�����E1;�և)��)ZȚ:!$:���&�|V@�) ���뭣�;%�|jB����Yu�Ļ+Wn�&a�u�mLix�|9�%���_��۵�X���$�Q�u�����VZ=v)�?�4Zy:C
O��rc��2%V11߀u�B���:��Ã���NH%�'�G�JǾ^���%��h���s�Y��F�]����tn>��c&׾O� x�L�}P���/8+崪t��)I1��^�饓x2՘��oσ&?*E�� �cw�%�^.���0�f|�y��@�8\1Ċ�H���M��nC�+�:�^\	�����_��ķ�i��m�lMhGV����8h���ݨg��!BT}t�؝f�E��5�s���k:��Rg�)g%�h~r�B�ha�|�˔8$V�$�G02�h�U�Y�b#��F�l�B�*a���3�c�w�1P�e� ;�� l�����|���z��}���%� N4X�uzA�0�G�8e���J
��8��$k�B�#�(����ed_�����da�Dt�����_��l�f[�d�Å-0 b���|i��j�� �n�X�p����u<`�_�E!�
/�Ѻ#�v��,K3�N^(�	�2����G<#j2o�{tچ)�?t���!�3���D~�ì&��"�&����-���K#���u��<󂌃�s��UQ�%k�~����R�G�\n��n�}�ВQ�)s�K�F����`��1��-�A[S�:�s���#w���ɜ�8K�%�诉�#��F��]�0�쏫8�o5�n���h��-�B�^�R�݀�%��.G��,�>���>^_�7RK�4��_�>�@ȕйp�Lǻ؈uu��U�i�)ecP�L��/g�'Y����44����ak���S���!6�r��
�U�/��B�����@�>��ni����⚐D�R��X����J�A�#�+�.�)�^�ߴ!SJ"1��W!�/����r�).�B� xҁB��<���E1��η��*s�F"��I�0G��z�B��(l��]  W~���[d&�N�W�#`�oɇ�S��y�*���#P�����޻R�
�2$�}��b9��WŶ���&$u)t>��vfi���8voh59�&=v�a�@Ee��
[�H;h1�"��>��W$��	�Rڤ�J�n��SX+xWI�ZP2�	�@BVB���22�B�ms��m�hkD8ρ"�1_�q]��G�2��ɰWT��AF��.,�Im֑��i�ͬ�s�Xo���K�v��ר�b���T�c����)�n�VWެ��G\�&�3�irȃ���?Oɲ��_��h��\��@����e0d��%!�e�23v����I2��v�<�L�u�<�7��7�)i9"����yԛ;6����0h]�)$����<�h��U�ǿ��xNCk��{�-2��*�W�e��*�L#c�  iM�Lt��ىu푖AM��"������T51qpl/5p��d]�ƥ-�˫��w���D:��S��UG�sU�aS�K�Uq���'�����;.�e��e=A��+6;�8I�Ʉ�C橊l�G8��re��j'(K���|�+y����5���q�-V���lQ=����$��Hl�e�j�-/�!�߰�9��j�ͭE<	oE-vۻ���0k�&�2��S��"��}85[$���{�D�$꼽�wk}�@Kid��;��D3Wg�+|dZHunG�9�vW�@�%z:�T F+��?�A��HA����/�����T�Q���+�~�]&�%������[�0�[������п!����?xи��ٱ�׷)j�+Ko��ox�{�g��oj�[�M߮{�}�U2�}�I�B��D\_�_����Y�����W:�p )P�2=i�O��ٞY�H2��^��͏ԛ��{ݝ+�۶q���Pw�lL��*�����TM6dX�V��GP����RY��h�r��L��ƔiL�,.o�o��ŧE{�iљ�����`x�W䗠�ʓ���?Va���dƑ�{�L�(�����a�^��x��guw;.�CQik�:�7cẃ�q+��*X[�V����iu�^,_���-*�� "�T�@euĎ"u�dGt�ʊci��$�{-ހ��b �8c�C�4|��0�8�7z��f���<ʈ���v�
�������p3��23���S3o��4(��Pt����h�6�j�q�r�.ߢ����Le��'h2�c
 }��Wm�\��վ��d���at�H¢LU	#�,�K~�krv ����$���U
����I�ݼ:�%��Q+��a�<�޽'µN?����K����ZN���<�J�Ԉn�?n ����M�S�F��Ŀ�rkr���+��c�޵	P$�M)��;j�c���f�&���OLR#Z��8/�JZ��=9��0��+a���>%~X��w_�L��݃;>Ơ�{m���^g���h��f����#��з��g���ΰ�p|5�L�=��?��p�����Z��2����k]�{1W�����V�r��v���#��
�{?wk5,Q��2j��\ ��kvZ����*��U�j-�<�7�~m�:4b�pg�ZQ�PoNe�l��gz#5�1�kf�����[�"5�0��r��p�a�^̹������Mj��#H�l!#eeyM �*�;7�#��Lj8�ю�lt�lYZ}�X;���_g9����l'��c"�QW$��x^چ)��T*�*j�������9\�\؍ef ;�f8���^F�H���'�������٫����9\�qL{�+�)��$���$i6�h%<b��e�%|��J�Ҽ����u$���|�ZD=$]V���^�>�{�:У��2��r�H��8~��P��o�M*��NO0���m�T|,*l�H|�� ���AA�	�8�Y�y��IY���oΖ�|  ~���s�`��잷�VCU!o]i�Ǥ������ākS��TT]fH�Y"�E��'�E?i�I4�r��&-�Je�i�CD���DlC�D�h�U�{�ˡ���Ŕ*���t�E <�+ͱá�:�9̼ �����=vf9���/_���X,����S6"9�Jy�$�?	��*�^�[˘:�N]w�8 ��ȿ>2c):��.8-)���ۚLPUB��.��-�ϕ��������;���;� QxZ�������5/���Pֽ+���Oc�i��'��o:��(�i4����5�F��,Tm�%�:u���VVi���q�N��L*��y��ݷ�J�21^�8���(���3�������Ð��/>�WF%?&�uNT&P���_��!�8�69�OxߐOky�F�`������!/���nja���%`�0���6����;�*���<|�Op,��A����_��3���F�4^ac�,	�(�8�ݖ#*f�"ʛs/��t]��.�X�Ҷ��Vߩ����y��	��G�W���[a;��"���K���?dzlV�n�[�ף�`s{'9X9:i�uS���!�N��JhA#�~ˍFX=��ԃx�[d��%;��q9r���*���j�IB��|���Wu�.��}m%N�m�k;2�p<Wx��G���$jtN;���a#!pNnux\tv��c	ר*���ߓ30�N|���@��r'��l�R�O��ﾔ;�W� ����+���T��v���J�`xp� c<hB�ܹ(=�S� ��k���
��l���?�׽2O�����$�ĲQ����!�i�(�u��d�B�Q���Q%�l�^�6���C�O�箈FO��Z�)�4��z��zk�?�TqH�uW�����A��DR@�,P�O�@�)�i��7�ͦY-y��Ҙ�ռ~0 ���v�1B޲�,�)�ٳ�5����jh�i�nC��Dd^����d4JƜ�8Q����"���4����h���-&~�Q5������1��~�)�2�t��K��d�#�P��
i�C9\Z1] p�l�,�d}��W��	c�X�7I�7�N]uL�nBx�纘?��χ�rG�j�Hr|�	���`��4a0c��z[C��z*�8��7Q�0����\�P���T�l�S�yV\�u)5Q��
M�4�p^�\^`�w�ԇ�|�j����-���YhUG������|���������,���@�؂���$#�����̍��.tA6�">���@�l��J����'X�g�V�J���{������=\�� kd	����˒t_�-!�6&{�[mHȯ������E�����29� ���P&H�]����������;�T�И�*rըG��Y������0E�6w]�q�80�C�j%�9j�quYQU펚ކ����5�v��aJ��x�W��ZdD�´�
]g�ͭ����X�O0P�-!.�s�B��,�#�댁`���;u��e�޹�ehα��1s�I-�g��F�IT$��q���(��&�!�[�.0���Gc��@�4y��e�㶂�G�@�rh�zS�����)��Me�_3mY��캾E���!E%��9ӥ���B�� �G~y�aaMv8�'i�q��1�9<�X�\��;��jA��* �Nm�c)oHU��0r�&��j�	��l����y�G�.�%�IG�r��rIT�
�5�'�&"҃���፠$^��6���3���c"Fy�/L9QJ3���	">0M�p�N>�-^9i<}��������G�p�!��L�x8�F��*�^|����/�`�zf<(�K	���b����
0"��-����-y��6�L��izY�5&E�m֙�E�ǙWљ���'~/yFA���8�*[ �0L�c1,w��5���aw�$��-|FY��%h��7�'oU��L5Qlx[�O�d����F��^	ZmъU/\9)�dt{��i�Q��۲���1����v�<��~R����g�H�w�A�K��<��t\:��,�}� G)V68e�N���:�M����+������-6&*�V�w�y�M��`���ׇڔ���-��+���r��.?�t9+W�����5r�6-CT���@~����q�[,������U���΅���!~�z$&q��v`6+������4o����$EG�gۜ;lOO��@&�hqs�	�1�����:�O�����R�z�5�G܉¿�����Qۡ�^T�����}�3?z�����F�?F�aV��d��e�B̊a]��m�
�U�"��(���ځ��*�W��� ��s.������)�� "�brX���M���V�؛�Ӳgx��B#��P�)�e��LtVs�8q��^C�ү�x�+
3������lW�ۊz���P�ϧ8��x���/��u(�l}u���*C�ڥ��!�k���ٜ�Z��K�+�u�n�Qb���������
����?�D�RHw,Y��B�ؤD𾬡������R:&�5#��x��Q.M2r���1H�������$��	e�-,6�.߹C�w����w
Ĵb�t���5�L$+�!�C��]	�}�����{P�f��1[}�#+[�O�����Cz$?'�(�Sۇ��d~W����$��\j�O��Y���%��1*���߅�Ŕ�p�t�^\�/I��J��"��&������������� ���tv�|�Z4�d';S��*8�g��W)����
�Ve|�l��#<.�*%�r����mR�D���~+��B)GB���Β
/.�<��ce�,߿�&�*n��>W\}���6�vI$���$:�CSk'@��f���F*#=9����Ec�
ek.w$���s_�ǻ�@��#�Vɥ~�C��z��+x �����D1��W�;�iZ��Q~?��!��[�y���NRO�<�h��ڜ��ۦ��%�գ�8�*�
	�b�.��"ţ;N����������{p|+C'�'�81���LI`�u�����&��F�e=9V�G)�p�p:e&"f�A��dŏ 9 n1�`��n��CFh�!��X�~�P�lNJ�ѤZ���@� ]�LG;��ц��B	�Ȱ��p�M��~�䄝>w���)%�M��M���S�a$�ͻ��:ο&ѕ(�kݠ����X�K�k�]�R"��M����y0C�a�Yг��G �X�1������W]���{���F��./�Ĉ~n��	�͹X#�	����kף�������=*�g5�`��Յ�azWD��6SY����!��F��љ�m���7�L��,S)>鞰���xq��_��kG:6y��C<�L.����F��'+��+���?��\���!b4��Ş����f�+
�,�X'����>���?%�攳�-}<�����4��+�C�-�k k7��8��y�EB�ZIz&��N&d ������	���q�q���|h����o	�M���n%��z�$�
h��P�";̵�x?[wm�~�^d�"��2���z}D���.ަ ��;�z�Np���hC3[���;Q�]����Pp$M�[�� ��m�1�V��\EcR-�n���U���
��i�B�kD�U���<��c��������Az��LS��<�gΏ%�2sU]ʙ	�륍SC�Y�0
���fL�V}���q�KLL����_@��hy�9Qm�"eYݩʣ�����`^����)4�	^y�6��jU*��e��L�u��-u�ܫd��:}�Cv_�uD�����ڰ%$���[�_�ѴRF��n2��m ��-�zg���\|0o��]������,�*�%If���;:I֗��K��^.��d��ȸ���7
�M������c]��,֔�Z$)�9ڰ�)��g�)"RAξ�M�OMT2\�r������[YH���V}��p����یL���}�	�4	�7�\��iJ�+�u�$
�D�����}���լ�̹o@�����"D>s;h�g�X����ҌP�2�{��)��] �pMp���n�c�ⶰt�V�Re`߳�r>��*�f��0�nn�L۹�}B@�x�a\��~
$]Z���j1��7�)��kP2���u�M�+т+J8�&�k���͢m1_2�G��ț�Zt1^D��f}kKY���t,��E<�C�i���HDt��+K���@��j�^S�Z��3ز��*�ݤg���T�9V3�ϡsB�7ov�,@9���L#�ۙ�m�h8�H����;2J�b�9�4|���S�v۶kܜ�O$��:��s��7�M1��G�	-�W�Gk�����w�q\�⏆�oU�H�`|��q��{�C�~�Ov3+q!�(�A���+����A*��P����&�_P��-K%�`'�p�6�~�\�2�k�_6��r�+`����.�/�:{ê�Cl�A(�֙���l��w�O�E�d���D�1q�J0'��m?��y	6������0J�G�^�u(�d�����P�~}��>S��T)W�)G��ء�y�żc��H�\�0����CHr�*;���+��^�B��(
���p�W5��.�[�9�~��{ Z�Q#!�b�~>�F��AD�����X'�j��^�HI��%����C�+�<	���\� )�+\Z##a�f�ϊ�xkd�k��0dr�Ɣ6f�Ug�zY��N�<Ք:K��-�/]L�&:Y��b^.B�x�]�`�s^B�^���ib_�l�He��!�6�]�`���}F��Kr� ���Ϛ4�a.�1�����w���<����P6C�1����6���5�(����a/u ��b~Ҷ��t�Qt�+$j���W�����.;�Ֆdv�'���%�)C
i��X�#�V����w,Ϩm�=V�"�T����.1��8�����j8*v:j���i�a|��ɵ]]u�bN��`
ѓA�GEVo�fV�+d�9�:O�V���&c\��F�bO��VE�i�:�SU�:�1��`�+��^�;�ZR:�)ȭ�X���T�CX.J��l�e,/�}��&4��17Y����J+5�3O4�� 6R���x�a�'����]�+����9'��UNҌ�S-́RS�f#W�T6$b��q�o��(��F����:���}��8կ����2T���D�a���K�'%F�,ձDyicѣ�3� ��
S�����0���;�yIZҘ��2,A��wD���̖�	\��d�`������Mz���n5.#��;�ζ\D�����>����Wd��L�pL�)�X@���D�P�9$�H�u�>t����vB�w+���� ׁO cM�7�T�j^�a�pX�\����_��-<ގI�I�AN��P���a�N�I�
�\��⻌9�XZ�b� /�I�"�]t�&Q�������?�a>�V�;.K9�R�럩������94����Qz���ae�� ��$��:Bc�	N�~zLH(�5���`�@8[�g�/.PFZ���7�B�2����2��Βū�8r�EP�Nk�)l '��4���T���}� �B��&����`e�ԼI��J]Rgf�&���?����b~��w�%|"r��(y�|���R�E$��><2��p�PM�a�V�m*e����-��a�C�A��lU:\�*�{�=F�ǝ�ǥa�_m<�:�I&O�L'�	�R�ӧs"�P�z��\�ipo��N/"�*�yW#sV����F�h��L��8'�{�UgDP�(u3vb�P=׍�~b�c)���u�{�C^�ŭ�]wE:nRz����AeX���}n��*���4@:��1_pZ��z�����F��8F��̤?�Z���F0L�������Ef|��}�p"���<}n�c]���h2SJ����4Y��Y���e��"��"��0�A쵠��c����Jn �\����?&�0)A�	T�UC�q�6�w��ս�jMzĩv�:�n�/�!��4��L�l�����oA��1�@Y�o�)�Y��[�40��N7ľI��4���_s6���9#:~P�hLDJ6�,���?]O�T�1{1��rqdGT2�/�J�A8/�3�`�`&�X�\͛�Qq����޲c~蛞|իT�h�r9z4aTi$볒)D��cp�VD�!���fK:A)-v�%Al��mԟ/y^	7�#��i�Zd�ч�,��� 'Z
D�e��")�fmmT�t��^�EI���p��������@����_�y�.��f��͋q5��K���� P*�4My�-��;��U��I���	H��@+��Q��֛�>��4��;A���O���&�������Q�֪2�3�n@P�
5��b�m��Il���3��Ϲ7�Sv�7Y������,g�pa�ۜ��q���:bu3�&C�_ڡy�M��}�����0���'�yy45��ǜ�ב�I�dḘ������$;�)��Gu������U��<w��٧ӒV�p�p���d��2/�����3}Ps�-PUA9^	#_�^�%b����8��� /Wjk��8�躖Qע�N�?h�������_�_���_���4ӽxd\���^�
!��f	M����A}5�4~�Ц&a|	��\~m� 2�Ydr�5u���$�T��Q��"�w�g#�d�/�mt,���*��aU ��59:�;�{8�3� v ��o�J�D����;.k�AM��t �m%��'E"�X&n�J��p����>3��m/ N=_Ʀ�+5F��ë���@T�ߡZu#�<i\J��.��C���"�5�}�T�w�#P?.�_�\�b�1o��,���k��w�q���բ����{�܁�c�tO�S5�p�����n� <�%aI&K=�ɰν�Y_����KM�k�}f��~��B�Y�.2���F Ie>W�/�Q.��ln�,�ܑ}1����ߡ����w���F���g�s�,��ᕌ?�`�
K ��.�ĩqW���On��C�hP��	9&B��y]l�C@����:N��u��V�7:�KV?�R�뒁|�^=�������6O����Jb{��aG�tn��FZ�|ؓ�j�b&���Ӌ�8�r�6�'U���׽�Hc� $�m��c�!A���躬�U��8��\iX �&kc)��k��t�WN���&��GKZ��<8mC#ۥ� �eUc0� �CG��>`��=���5�w�c��Έ�5_���J�7�C���Eߙ�zA�:�� k�pa�Z͋J��+�+f�!:��^��](uZ�OvdP�E8��}[�4�P����_�e=,=BjKa]�9��f�PїZ�
���)L
�IS����fp�t��H���yH�V �� �W��J?]p�(���֌��>�a���J�o����a�?�I��v�Ѓ:�.8���8vx�8�Gx�Gͽ���KQ���l�\�G9���g���&��V�� �C�C�/���.�P��='$�i��%d�[�6��T3$�2ם�wi������~1![�>�ݢ�Αa{|i�h]�MF
��)x��6�c��k�ęc��c���o���}��n���
��|S���z�ѕ�5}�wJ���yw�a�u�FF���r���]����z�Q�>�E3����b��E�C���l�n��t��b3����7���1����:�Os�"M=7v	��)�q��_�"#�bj�����M�"����,��_��K�+�5�#9�zr��|�n�/��fy�g�p[��ͼ��'J��!r�[8��sAʊ%�~bBe6Cj1=�נ��ST���}a<��7�|!�~U��Ǜ��&�`X��_NJ
%v A?=��'��+x�����M��Pz��4�:*�ҫ���u�HA���0�V�����r(l�����o�ã�snp���Kk���7����P��Q�����E�>���[�T-�/-M�%Ԩ�aJ���t�%�7�J:_b��dG@F��-�F���}���.V�SY�(S9�b/��C������][�C���o`�Mn9�6jk�F���"�)�Ξ��/��@#;�)r���uł]y7��s>{.����ve�b����	���6��M�kF��x�Z�	M�@����8�xY��f��o�;~#��!2���h�M��EcC������&���S��]�<��tǮBz��w�\}v`��>����`�⠮�{�8��H!=�C�*�|��F9�n;�����������'!}��a�/ݾC�Hg��i��;yaNW����l��Klr/AW�-���u=����A`��ʎ�1��֊�R�JZ���Nn ��$�;Z."�������4lr�֋�5�8tZ(��������'�y�[VD��f����v��]�5��}F	Y��M�'x\Ǆ�1z�
�����
z�B�~t<���OW.���u��sd5�b��)a�D���7ۇ��GD/�{�%������_w�HH'S/B�2�����?��1x�в*�l�:�A��S�pw���Ga)�,!��!�FC��� �gC�%�1����8X9
����KU�V�e�R�<�?F�b����;��a�{t����Ä&�/���<��#(��Zx��
(��J�#d�^�^M2��ªO�钿�=ky���0N��G�t�YO�=ܒr�`բ��08 �[���XD��<F���s4�'�@�64�W���>���jإ���V��d������Zc�5��RM�cv���$ޠ��:��X�j��*؋��z�.��*.fQ-��b�}z�C15�Z�GT 0ĥ$-�}�����bڀ�|�k3�濭����(��We�i����AKv��<v��?9Z7�9�P��-O8�S��]�D6~���p�$`d��.�$b��X�R�Z��n5�۠��M�WŖ�43�[Ԕ6�
lrk\��QifJj�'��\�D�K0v��k��x�n���{L�~�o洡�t����x����HÅ� s���3w�;��Fb�ݦ�|��sVC���+�9�D���-�v�֎yAo��f���)����Ro^Ƣ9u�L���)��$>/Y����b� 88�9�?X��Q{2�q��l\Wp�R��XN��)�y�Z"S^"�0���J�i��f�m*-p8"�J)V��Qw�)�2kO6��wB�#k.���s�dl�������Ւ�ז�h��D��u1V%�?>IhT��r;:*�̲p�)a�?C���7�yKh�^�E�rZ��mG��)B��A�� ��ǍI���#�(�̀,�XU�8��4�!��G`�?��PA/�D`�����V���;�ɼ%�c��O�I��u���v��6�C񲃽�֤C\�hwu����l3Z��>���%�W ���v��	�YL�5�mx���A���n�6K�aF�иGڄ��fq|6�u��%Q�H)ۆu��P�� �Q�i�װo���H5�7�i�Yv7��B~i�� Iy�`���~0�L�20J��3�w�x��y�Vm�
Ă��K>��(z��j�`�}���9�����`] ���% �kr���w�W��BuҺ3�N䯲hb���n�m{�YAOM#j�}�v(Q�������-]PT�h}���M��T�B�M &���>�vk$|
���rT�\�\?��̺[
�?3X!��8K�^�X�l�;m���C΁_c��E�^j��'��Iz�U8�ܺ��'r$�ԊC�������x��O�9>������&�ֺL�ȣB<��'���й���J�=��˺�䲏+�7��� �s�	�<�̳�[G��e^$VH�S'\a-�zܔ�Po/�JD|�t��Z��l9��#bq���<:G�Ps�K6B�vj�g`l�}�5MF|���Zz�H ,2,C�xz	@�@����Ց���Q�1���1�_j!9��UCq�[9��eRUVhe��@���
�ʅ����G��	��_��E�(������9����!F����HNv��Hi��f��<|٣�s7�����?z����Dl�Ґ#�r�a�e�FA<*�{��w�w����e���F;5�⢢�&���<���F_��ı�1L�S�C�>ar�4B�iz��p�Ψ�y,v�r�,"�B����<욧rKZ\���;���� Jl}Wy��˂�r��b߾�_X�*1�u�%�x�Ķ$EBi3�����$f�	zf]�T6�-�xx9��� �H$/���L����O�Ia��OS��p;���3I;n�����O{��8t#�pgB<ުwn���@b���{����?��w��+:8N~KJ��V�\1E�
��8����V��7�e�lV��$�_`3��l�a�&���0�����ɮ�_F�`��ȉH���yTOz+�C���/��E�I%Z:�_�Ob�dR4~KD��>��_\:�
�:lF��򹓔ъћuh:a�4�M�<8��"��>®d	��+�q�z{��k&�lTx�����3���]᧌cUV����͟3�գ��1��R?�0��y�D��M%�Z�k*��v�!׍�X�(�[??�4+�;l���B$d0�hB��xAq��:�0�S[X�"�$�Vڃ�	y���S�c�Jn����^�NtPX��rڣ��g��'�}Aǂ�!�.�^D�34�ĭ���~������b�O3mde9�p�Әq�	?���y��K��?��6�l������+T�$F4@���-�!�� TL�zq9����)ͺ5�r����i3;�E��Fz��B��=b��lA����Jm�u�L�*C6�l��ط^��wUџ����mc5��vY���Z����܁i�D`�@���N�����	� ��-n�2F�6�������0����ɀU&lE���Ĩ��>Żs��h���z��x3�D$Ĵ,���h��Bc�tA*F��m��l��oI�/$YJ�^!T�g������;��]u���Ɍw5B3Q��O!�9"_�P�Oh���3�(t�[�Cw����J�Ϩ ��4�N�A���1��u*>�~�-����t���� T>�:������I`-�tH�a�L�j{()�'m+�Y{pr��>�	���i>ч�m^�*[���\a��ׁ�l*lN�1ɗ��\]$;��:��Τ��N�Z��C�Ff�zH�*WlQ8W.�m+�X���+܎�dL�V��Rz="<��;y| [?�=AEg����hc���#����ݤĘu�_y�J�\���f" fao*����3�+� Y���+���p'���Y��W+_�e�lo�d�O֮u�ҍ���Z�ZT?t<�V�UتW�ϵ�*צ�g�ٶcd��y
��˹�,�G[ґ儇ý[RK�s�����⢚�;�@�|�A"�p^n��v��U���clV�����RQR��F����_`r�`��(���ǫ[2{�]#�L��6�YY]V���8rc1���N�-8#o:
]��sO�B�����:$���#di�`���XGǘ�ϑD ��wS����r�߃;��SuЙw�¨K�*�`SR!�ac��E�G�x����Ry��ҟ��� ���!~��^˄|s�NM� M�H�FF�=�����N=������QuW���߀�Q�lð�N,z5�c����,�&��UL�~�f�W� ��PFߘY�a��!qKRq�
㧞;Ӱ�Z�
:�R�jN��� ���G�{�3�#���Ꮀ'?�����33��[y�V@f?��,Rj�?��s����$g�r�;��̀�C�2i���s--?l\����O�-u��:[&?�UH���*�y�f�V4�.�ŷ�d/#)�e���b'�'�(���y���v�0�!�A�`{�4de'��/v��G���C�@dh ���*�ޒ4l
xh����x�a�*��Y*{4q?��W�JMP�Fn����y��U����C�%w��)ټ(.�.��Z�d�/%�\z��uel�`��s��C6��6K�5������}͡c�]���`��,�t�ݙ�rΌ9�z��6�tF�Ϩ/=�����V2K�'�ֺ�4T�t	Pr�ȶ4�{�{�%i7����L����p~���8�\�85�ڽ�k�)��S)[����T\2d ����C�g�;�4.��NWީ"�b�%(���+�t7���CI?PMR�	�ӧ/c����+�^�[�29M5�Ւ*B�r�`��(W�����Td��MdR�i���Gm��nʷS7����	Xz�IJu���w�����ǈ8V$����u6�]n��=��0U���WX��ۤ��'x�l=U�?��u��%R4�(WB��(!��m��[eN���{Jz��a�U]CW�� �UTd�K�����8�6�Ї�!�	��G��tgG��{)=�d�"�=]�֘�¼k�G���i��C`h�?k���=@��$O7�x|~F¼��!$gs�F�:1Oۗ�X̪�WN	�f�f6�Ӥ�gM�= ޿��H���G�#V�2�����P� q<F�^��;���~�^rt�=A�)�݊������#�G��p`&>X��"�:���C���
�S7���C,R	Z�d�U%�.eB�O�l�J�L���t�Q^5.�A�Ԥ4~�Ya�fѤ�$����6$FJښ4D&�0
L�a���>��lѼ�������b~��Sh��C�;�:���
�꺇n�L����l�^6�?�����Q ��vy@��/���-%�lYhZ��x����j��*R�W���f��B�g8��N$+�ӭFP�5֟���\��s����"%R�j	�N�B���͵���Hݐz@�m>:�C�`7���M�#v-,�d\�����:߬�#��P�A�s��wh*����|�2;ٽ�V'��6��q��$�y�}x��?s��Ep��5�ɭ�,K8�@0��O��q�L?�o�%�3��8&և���xvR��5��tG���/�>�����ofc�H�1-˱��iBx	d����J������#��J�}��*͔[�o(GΌ�5�@�f^��g/J⥒�U]��46BF�q��7s�mz4c�i�����»x�}ص��x���sm�#��#9a{cbU2ȡ�iOq���Ϟ�c�Ƣ_#@��nK��\�Eo�3��L���zB��KM�e.�u����ɤ'c���5Xr<�M����+�H;J�B`������خ�_v��dW ?�h�e�Cմ5��@C�cx�>��&����lax�nu+V�r������Nց���<��Je{;M�0��������sA����Gc#=N�'w�}~��j"��]z�������^'Ky�]�WR�����Q�s��3�X�n�0Pr�"C|S@����`�� #J5iȠ�r�m(��>	E{XH| /�-�w'G<	���%R1�,�P�*��r4��S�o��[${��=Q��09P~	kf%�2��׏~�fc�\�x��B�8����Z ���H���SEp�D`��O�m���nnQ�S�+�+�j���#7���Ό�f����ܩ �M1�I����U�z3��-<}'m̲**'�����d��~�6��V�!kn�`��U��j�lF���տN�U���6�g�8p�!�٢}��W���	�(����v�l��O/��27g&��Q<�`�!C�j��ӌ}B!�����j�ɍK���M�5R۳$a��QQ���'?	�k�����9Ѱ�\�r���� (���I'4���ٌS���䢺؇�l���W�(PC�`�qO�"#q߸��~�]^TtZtqj3�`V��3��q��L43��.�/�K�B���Z9=�z~��t�[lM���Ι0��e':�en��w�2,����k*�	35M�<��I��(	��5�1�j<�qA���N�*�f0�3�B�{�J� *�Mou������bG��N��̜cc�-n9�1Q���+�h����0��z��ϥ̋�t~mC@�]NDrN�a�|u@p�"Z��I��5�!�&��X�hÁ8
W� ���!��o�����骸`�##4ڦ�a��+�ϜF�� ���"�Kt1�F��]�Q#��yۊB[�A(���~gMΫ`�r 	�ʸp��$~�p~���-������<n��
������×
f�;q7����D�	5�ξ������<3 [}Ug]H۬
n��X:�C����q�x�/�*m3��vS;���9l��Y�	$��i��M�4�tC>)l�G;+\}e��QW�4�m*�n:d�����r� �5�?��Ap�Ot�N;�n;��FxI;,�f��' �4Nl��FdR�
�gx���a����*ƪ]�=���1sc9��(�--�4s�F�G.K.U����~��3.�=gQŢ	�c�"��W���~�0�f
�g,��Z��`F��7�6�7q�#F| �9�b>T�������Ǵ�,�0��w(��`��[?����N�J'j��UX>t����.����UJSii�ټ�Xˀ��������1B�W����b�F
�d�p�(7(RX� % �!�%����_���ʣ����X�P�M����ÞT���"΂�Pn~��M�n�Gu(�|���;�+wk�.�Ar�m9�^]'u L)�qAx߯��9��z.zg�}��a�# �Ś���.�5�O*W��z�������x����ְ�Uʭ�������+���.��$�6�Ю��A�+�*���+9�$��[����=�Z�5��
��ĲЦlOakQ�B;]��z�>��ۀ��lPO>˅��@��`�p�^� d~����m���Q}L�)�"[,�Edv�y�<�`R��9AI코�3V/�����-��>�X�.r�	���g����U��_�q�,߇D�xwZ2n ���<��[\������:5��^̧ȻU-'�=X>��+1t�ie$�_�r��?�oBI�_� ��ۈl%_����b�'I�j�u�l��/�nqO�-U����,\��������.U�_���|	�v�l�B��c�]6��3��C�a,sY9�� �O��87���EO��狐os7ʭްZ��$�w�~��CZ3n��U�^�<"�Ǉ����'���a�}�#����O7���G������ȷv�"�Ի0��f�f��i@�=Riy؇Æf��tRb���je����{鰒�c��X\$Bȴ� ��ˠ�V��v)"4��ΎQ�D�V-W�G��-ֲ��q�]���J�8ԭ5���,)�Řq"��������Фr�D4����{�Pީ9ſy�tCr>��3���a�����8�����q��UL������y�0��N�\��t�0�w��WϨ���9���)�_����S
��NyB�&U{��8�w��*���w�~�J�Q5��:X�M$�\*j1V�n,z>@�� �h�h���2W�=�( .tc�[>"*�j�@��Cls�bG�H8��r&i͋8�P��kU�|`�R:GU�6�s�X{�`��62�e�>�oSy�)�q�cXJ9<��E��!����s<�0�6�xo��#�A�!���$���.7�����Z����\�s�>e�����wp�O8������r.��%cc2#e�]>���q�2H�c����r'��OF&��ZE�&���w0[�T���5�>�C��wZ���R��<�?^�����ӐW�>	��U &�n�!#rw�l	hRbS�q�(v�p�#x���ሴ��˰�[��(���3Vw	���wc��d����ֹ�p3~�3'3MԈ�Pr�~p�{�����kg���2^���]���[tc8�؇�Jf��a��&7Q
(�ov� �LuSޭ	�}�3� �'����e�n�R�H���!�Xg��d�u-�Fb0}b�~��	��8�ş�U��6`FU����'�rZ+ځ.���{�a�'�#m�H1l�n�D������.�/��K��ϲb�	���:�ԋ�s���Q*��0�F �}Ď��(�0�x*t���(Vذ	t�!��y'w�l�����;9����e�O-�7�.-U���G���ّȖ�%m�LrdJG(��#j��� �X�Fh��������\ߣ%AȠ �j!����s�<��ڬY�Oއ)D����A�u�95_a��PۢI47w�=�v<��u�s�5<��`CS��+>,W���I^����j�֊<�8@:��e�B�!��Y/�?Cy� ��b��v�/��km`���$;7���e���¡�������	����|��9�v�p6�~
�xm��GJ%��؊����[�S��<{�Ķ���^i��X���QM�f�FT�k�i�/ZFQ�Q�u�u��VQI����
���UMХ�1�{����c��1�Z���'|��� �>X�tx�>beO;�b(;�#��@�4c{��x��6H�_����%Xs�Mʨ�n�QQ�C2Ƙ�I����T�2u�5���LS�%ޓ�/����|ȷ��`�/�ݏ���<Y=��0�V�%�����1n�.�G�Q)�ច��Ɗ74��ć{��������Η+u�����	�N��kl�g�e��C����&�^WB���P����(!�J��W�-Ծ�%O`&��e�p46w-����?�@�R��EC�wU������\S:\}�>l������l�L�_�����^�$;z�&>0�iHܠx�(�%	�[Tr_��.��t]�G.����A|��x�WL�f�ၡfF���<&\
�q�:RH���˧A�m�PA�������Ukc�g&*^'j`�'��eFaq��݊��L�)��$�`�0���n�<����/��U/�>`��#�LJb���U�w��n���].dNaʯ�,�էE���c\z,��( B�N ڋA+���Pz�:aӯ���x�;O_,���D��ze�f�C�zO��B�i�ؗ�e�w(�=6C��!ǒ2�߿��թ��jX�;��m�x�_�����s҆���F�u]���ܺK�L%k���j` 7���4��Hsow�p�V,��Ϟ�J�� b�ã�ojΟ�N-#�\��`5Q�z!�u��x+�� 	#g��a�wo*�^Z#�tjmHl��[�GN~jOw�r`Ю�LPj��e
��\�S���4��G��>?�)B�w��:��@y��93��� ��@�vͣ�Rrj�g=	dW=L�5�G���5~�"��2���]>��u��)�y�b�o��/'����
m;����O�|��<�"���F<�Ok���&�SO��
�r)�p����->�����	��jM����+�����8*bOl�2;:������t���B�OӜ�G�~V>�H`��/��%���D'�Ѫ�ڰOa�V�+G�%��@�Dؚl�C��s�R����[ER�oOli�#�_��ȺA]ñ*�ꆳ7�ƙ�v{�ޅi}���b�
���K�|�|��@@	1ٻ��E��l���@�0&��t��'~�	"��wh6��LYy}�`X(��`s�^��o�)�K ��M��Wd}��Q�L��E��K��2s�2��:�,�pT(�/���P7SeZ)sF�R2���G�r�rQ�<���W�n$��[�a��WLle �P��4�`�7�<.��
�>z{���cR~ix��w^�oUG��U���~̫w>a%�<!wk'=v��M/+�D�(s�mf��{�l�1i�4V�k̍dJ7��J��(�ɯ&��(�7bI��n	���\��	��x�ks��l�vg$�� ޲�����I�U����R0�Z��nFۥz�f�s��`V�&���Io���T��A#���M����1�����z�b�6O�[-(1�،՗�V��Q��ʐ���R�p-B0>Wgˌ�E�Okw`)B��Ue�	�j7݈`s�3W���8���� g��_p0�:�u$r6n�\�tPH��&��eWh��x���96�a�։���Pe�IK�6Oh%�-f���D��v3ב>DԶ��G]����^�<�<�^���.��ߝg*���-���_	ӃQ����$x��#G��4_U�,4�p���U!��m]����t	2�Ǹ|n�R��H�����m������O��k�,f$��c�����Â�O!�,�����JC��uu��U�h���?�0#��-�80���yC�Ʌ=J���2��uHކ�
aP�̀���'ެ��sK>�p,��:.,h�}#?J/ro���P�<�;q� ����.�x��� ��_���TK-�I�m�f�Q� 9ikc�󌖟��j�g�����e-͏��B��V�U�*E�ڋ jZf]�E�q�t.�%g�F�β�wW���p}�T�\���Mѡ�/���a�t����m��%��F��;9%|ɦ�M��y�~V$?�Y�X�Tx�r0^��1���݌�� 1�]Ú����I�"������y�)@�����DS��O���'�/�p�%�%�n?Uk�guN�B@��X8GJ][���I�����B�m��������#�ӖX(���n�~�ܠP<\�Us�ڍ�';��d��i 8T�5�SY�ZYW(hl��k�{/S2c��9g\ag�'��6k�#�Tm�`ܪ@��FרT{XX]儭��-U�Ӧȵ}�Ѧ�Y�f���N�ӛ���x�L銼F�0cUux��o'�����_����s��@x������}��B]�C����t_���1����[v�$ބ��4�·��Re�#%1�l��!�+X#�G���X�	"�d�7��A��oָ�΀�.
�^<�~k����
�Q"A����#�Ӥ��V�vR8�Y���_���-9�珷=�u�eP�g�d��a2ι��3�
����#͔�� ���H��%����M��#�,��8\�h�����Z��%%��C�6T%�C��T���ag�on"��-r��-ӆr�����Jc���-��!��4��� ��@p�����d+���p1�RQ��]��8��-sV@rӬn�hU�O�5&=iG?i��~��6OWڮ�fUtK��>��X[,���M6|���@��P��j�OT�pjOkJ#�A����\Bp�N߯�uzm�H��w�0��j�������m9N��M��D�9�Y���Ce͔ڻ������q���"���נc1�X�aC׿�=�ae"S|~��,����0��l�|�(>ΠIP��<����7��7�ݰ�~�*�w<��F�?X���r�	���JQ1��Ǐ��z��/tP�u�zor�K��j��B0Bl�ʯ�1��S�M�3]��!��Y�bx+�/:�1�kA�����W��X����E�~4y;iP� ��FG;:0B�N���hb�u�����;�ֿQ���|�-����%�Eoo߀�o'�}�۸�����XT�rU���)�@���:(d���,��2wc��3��h{uWP�bz?#z$�s&ab)�ǧj��) �H�z���� �|c�K���`�0y?�0���ފ/��+��
Z	�U��?��r.u�4/��؁�z�d�;*֝���s%0@K ����7��Q��o�;Xg��WEڊ��ֶ�@�i���Ę
�O�4��`Y��U�l\�m�{8�]TG��ղˢ�3�b������K�A��E$���Wh���qJ]�ޠ��^x�p�s�>e@�9x�3����$��sV����kdW��\qړ�SQ���A'ni2�?I�1��:��Q��=�f��&�a�3ߩ�R}�+�~O��r5�_��� %n9�N��1�Xzm�}ٱ�z>��~��wY�6���g0j0>�$�l�	�7I�S�}Zt�V����M�oU[�u�"ѢS�j��)���Zd��O"u������e-=#D�)�	I��E���u�z��k���U���8#�!�I+T�u6V�kx�ܜ\+c>[=/����~Ҍ�1/�:�����&��#
iH0D#�	4_^/\�������S>ђ��n�iwX�;�lf���*@��rT�6�ZzB
�Y�*���-�
�2�]b��3�ߋ67�@�u>���Ӻf����C����~��L����kX��.���%]hb��^� ������,
�Z�0�y]O�Jy^�S��<�w��Z?�g�_<P��Y!�Lf此s�.��Wb�B�*\�,a݅Nr�A��p-�nA�_���ˎƖ���[0G��5A�A~�L=�qVE^D՗H�JaMv��X��ZR`}}+V|�����ʢ�3�$�Y���W��=�����4�_��x�x&�� ޝ|���S7�)3#��ͫ�S�	�(2c:��&���u���~���MP��f.<��9N�����)�M0%�O\���v8��KJ����%��V����ǟ��J��m�8ʼ܂�ϕa�����y��Hv\ry�x ǝ�8g�-W+��3.���W�k���I��~T�ZT�Q��5L�P�/z&�\\�)�F�����H�#?�4��/=w�
Z3s1͊q�#��2f�{��c��������(��	��W���Pf�|�#�V��A(��4BE֌(��~>K��(:�섲()QW�s�/�����������=.��6����j��	�����{�A(�#YO�Oݨ��fF���mJ��S�"W��)�R���@{Ty�w��m#S����)����{^с�&U��\�t}7/�~V=���Ey�b�AȄ"@|��� SSQ�bSo�~�"��L��A\�����a��@��\0�b׷
�B�HU�eJ�����W�5G\<W5����qF9f��HqC��E�-����(�@�l̔��I�(���~5ΰ��v*Q_��uѸZ��#����ܖI9����d��=Pq�fK.��8��<{I�1��'ȩ���ޡ5�)��.O|]<��A���}�R��]�
�|(z�$���sl3?$�R����2�c��*v�?������2�N�w[_�YI��|i3��6�M}@���o�4�k�@��U�cqu�:��iX �r�����!+v���G��W�G~�8ܺ�X����Wx���VS����O�f��`�$==Y�C]�4j��O�xV��3l�?_��(2�%�:''ݛ�s�F�74��'�!�0��,��U�aA�ܸ�d.��*��O�U@�a�̪ٗ��"R3�nN1�EO@w��Z�ഷ_+��s��iOUv�F��o$���G���ڈ�1{���%E�.Z��*b����~*�,Wl�T#<q�"E�����"_'v�։(���~���D0B��!S�Fr0mgV[k�Y&�G!i�@n��)�	��T�OǎԳ�����c�>^h�B�Z�<�~2,
���F<$�F� �d�ӝn���;�s���_�7���ۡ�t��O�\b��K)��dz�3x"� %��6J/�u�!ײ��k�wL���)��~X5��9�W��H�NF����#�:cV���T�x,�� �8�g�8h��Rqֈ�c��C���j�ff+��.�m?��]�s�&?�`L؎~���w���`�%���9ma�s����1�iv8 ^ohuvm��zs<�~^W��dQ�:�:�>=�>�$Θ�nى]?�$j7���h\��r���~y80CTΨ�1e�$(<�6tCJ��몦/�ݡ 47÷�Z��B�|���oh�8��_G&�Б�'�g��P���Nl��#A��i���/�7�e�-�|`�_�`�eޫ���R��F�f��Dqɏ��"�����CH#p������d��Q��9+3�Xe=�M��*qi���t��B@��-�=���0�դޚ�#B���n�|D�ü���f�qN�Ʋ��ݖ�m+М�n�
��{��h-h�~�6g�h��x�f~\�'�Ͳ����`tvq����)�c�"al9P0N�%#�Ć�ĚDjPk3E�R�%݋���[2�Ac�A�ydX�\Y7����.3t1@��?1� ��g�Ri$���M��L�k�XO\iu�j�e���gF뻠@�u��P�d/ݠ���#�� �n�����O�w��m�PQ��^3�K�Itv�mQL�� ��&
���#���ݦQ�
YS��A6:+�lS���#�q��p@(�en�:��m5��g��a�� <�+��q4�+��kZ"���w�!����F��y�0��H/�6r>��C0�KM�iԂ�SV}�	��:S��UO�u�{����p��1�j��Г�cEa����*!G�n:�τ����y�ߌ	�nq���J��vbjxT9���,�^�Ľ����V���CLz�˛_��Dq��par�<�BT���L8�u(���>� �{����\��ǭ�f���Ј���D|�m��OgRGFP����=0��pN4�����܈�t��:+��x'��!%TQ2#��4�m}�A0�2K�z<#�d�LTu�#d��"�+�*��"c��~�C�¨7�HV˝ٗ��=�1�f�yƋ�����Uٛ��P�l.h�W֑{�5:�̼'�j�(RF�����NE,!A9%�3$�v*\�}4���o�A��^W���M�_�y塶K�}J�[s$��W�_�����?��=�<.WQ��!�OC���~��c���%YU>yh����r�t���Ң��4�]�9Q��$2�� �9�Q��F9�T-ͯȘ�:m�w
�i��x����Ǯ����^�\���#_�գ�'~+}��¢H=����K��ŪV���I��O�&ϭ}v�A�����^��Q�o'Fՙ��&�-mEܴM��Dd�!X�����w���?���������:�_�_,m��06�����r9/c:��V��F`�5X	0)IjT��L��?e���E-�t.r����17�4V��6�%_�[̦���ӏ�9_���'n�\b'c�����I��gq �篂���$8�됴��)E0��l���w�+B��T�~5m�����5�`��}�o���ԃA��o� �&�T	�k�H�
�+쁐��r'��t���hZ�x2���[`��h����(�i�5z�[�V	��3E������Rػ�/E���t�]㺽h`;�V"2��T{S#]��G@7�+�����k��o���$m�~z^.W	I3j�9��"�a�k�cg�f���š~�K�*2�K����q/J��
nl)�N�
�#�N�Z\?��{���]��A����'��m!S���5d�c|��nwBLBƊ��7��� �wd�p롡�zx1������%����E������a����< ���F����Uȧ�oʏs֛�_�m��6x�<�R��^�7y�� ?^�?����B}�ls@U�$ޗc^YR�����iT�?#�z�H�d�=Wa�Ꞅe��'�~�}�xW�.����+�v�]*+�&z���ԁ��4�h�o.z�v�	�ᅰ�!�����h��9-�>�*�
#��Ep��E�4��>[���sE�l@O��������R�bb�	}��Y���y�<��2�C Ԋﰠ�;ťY����΍>78aY�q�pE�R��a4\/{!V��8R�Xx6���ҧ�P��`��8J1룘��򕭘*t�^����p�)5Y��� ��4�>�@�&KN9P<F�j7O�F6I0*�,8��f��{ɕ�Ʊ���I?�$ �zdp��s?
㬨;520���!ivq��+yU�a}I�����`5��l�<MT�˥䖂>�K������+��	��Q�P�9x���|����&90J�P ����6��#�%A��[�k�E�U�FC)(��zlY*+��h��{�e��}X�=�]1Ky�ӡ=}dj�_8;�aa;�=�i6�}=�����%��^�����|�(�۠n'���ɁH�Qϰdᣯ�c ϯe��Ά�S}�<��I$w��a�;E'|x.[�/�%;�=�����ߩ6@~'�"��;�����z <Qf�l���[-W��W^��V_f$?+\���W��aw�H�fc����\T�!�²�#���z�i�������(�����]���j�(�ļ=IP!�T��3K��	�#�{���O�NW�;ԿJe�z�J�G��J��_|�4�s���l^��{�y&�nc5�Oӕ�[�W���Ig�2�G��F�ӑ�2RҞ�؋��i�I-)�=$�<M3�|��_B�����2�R լ��>�<��П���hL��v���B�r�ҭ���)"p7	K�D+��,/���'	�wa�	�$j�,}���!E=����-�l��}�Gٍ���3r���L�bvw�u��b�.xc$�g��2y�6r��O��ȕ��Ӽ��v������Ԣ��|�nh�M���ߖ�sX�ⸯ��:�<���2-�υ�]ҵ&E�,D>(���E�^"+8�X���z�͉Jj���a�� +�,�t$�i��z(>�ΰ�� ����T'�]��,,qɊ������bo�>�{�7L-��
YZ��Lj���;Pa�W �c��ds?����W6�V���W8a��E�m��9p�Y�B����]<3tF`g�>M��/�47��}W�AZ��B�6١�8U2���BS&������ޤI�#do%��V��9��`[>�s�x3�6ęf��|�,^�����
���e2" odPn��)�%+�՟ ��̕{���pv�@v��z%��
��'͵dkm9��^Dp)���7�䷿��j������Zjl��2�`�4K~&_�0=�n Ez��C3��Q�
�8G�x�uR	@گYor�*�,HS__�3窯@������Ҙ���lE�t���	5��|��D�O���Rn�ӂ�_`a�/�7Į����m���O�Ǜ�ڠ�=d��&i�w����c0g��.�H����C(�jg[L�C��.m���?�o{"�sV7�_�r{A��k����.&zMĥ����w�K�[%XϽ���go�۬�Q��9�F/�:~����T\]��j���r����i�	 L�����	�<@3��%w����U�;���b'sg����0���C�	�ý�/t���M]�QyF�o��&�ݽ�zL7�B>���*��Nh`��z��#.������Q�������I�lH�h�.s3��X5��҉Ѡ*s�i�p���=;��i�sj�:#`�|���W � ~����uY,�&oZv�����4�PӁ|�>�@�Ɠt ��W������3�R��WjdQ����CT�T�����{B�m=�,���&���kE��po�i l�m��7c�\���.�$p@7�%���^5
;�J�U�'�t�\�VQ���{�^��;��S�(�������&�RL�S`�B
4�ó *zf"y�(�Z�e�t�mc}<����[�US���EAB,�!S�E�&XXA:Tn�sƃ�ܑ�ZbWN����ڠ���s�KH�k���S~�!��N�&0�c��V��܄�z���0�t΃~�-�2�x�o<X��MHV����Hlh�/BnD�[i���!�5�E��SlC��p��+���歏[0��_:B+m�&A��o�hck4�t���1|2�b����m�����4� 0�5U��e��%2R�
l�ʨ��et1J��r���"/���"L e_��V���c˒E�?qx*/���hٝi��Ɇ~�/���UN���_(0����l���8����d�ms�%�_����Xu���+`Ƨ���+|�N���������R{�ߴ�@�<A��rO�s����d��e��`�l�k�es�`���y4���d�P,�;ľY�������3�IJSFh'���~u��"�`	��$F��(SW�b�%��:�X��P��7V�*B�Dw������ߚ��"�[S�3�[�ν�1�5	5ar|��24⠈́u6CD����sdK��(8�����7F���vC���ʞ~�+~���D\�3�ouI�/l��b*�/EB�M��Uޏ���j=�v|B�% �i�����X g�ǈG��D��off��a���B�C�2�Ef����;i�|�x���F�+���A����/�C������9D�o8)�����+,Rdd��Ec���Ӹ�/b4^\I�>7��@��ۓ��*�`�h~2e�"�/.�U��"fp���#�aT<�j��:����רi�\#}�fq!^#�Q�����j�:7��0.c41��|�ӥ��&�`e�y(�'t�8|� �7��<�ץ:+l)�G���'����M�{������bA? �W��S����/�øe�n�[5�v���BΩm�1�Ir������/���+M�nMK�Ka�s)�&�Q�M��\O���XmI�!ɩy���:&&���0X�S�VeѠ.�6n/��y�C�y�9�Rt�^_��W|E��'=]'ܨ�o>n�+?	ԶM�Y7��M[�1q�"��� eD��d����Ӷ�0Y����\4*���@�*�)�n
��d�D2�]��A�8�M��~@l��7m�;�N1VxT�����
��LY��B�D�er c��7�����ǆ��n�����@fJGcc
�e�I�@�뼜1�9���ǅ��g�"ڤ��oZ���ޛί*���˦,�`|]��@�V��u���@sN�?,`i�4=,A�t�f3#D�f��t/������l%�/�-.)��c������ڪ������Hm�g�i��&�t���O
�v3�$a�x�uB+%�C�|L���4[��t�uM���g�m���~UX���/d���#8���t*�)�=�@K��p���e��^�gQ�j/�K�b�]�` ��#Ym �w����v��;��G2��x�9�g>��]���Ǭ�\l�W����vw,��z�hɗ��m�c<����(+�}n���������L_�w�Y)8��
��<�'�����}��Vɇs;��xB��a�����&ӽ�k(�on�`����Q�-��Ұ}T|� ��[��k+Ȓ��2U1��j+[�,�ɡ?�!�M����]ϫ��b��!$�����[���>���sv'<�&�%k��K〵P}��c)9]v���Vw��r���|2��@���'�:��}ґEqFw��= ]���(�s˟X������pHeIel�كN���"�:*R��KS,���Zc���]Q�o�u�����c"&*������(��'�)o�?�4�L�a�&�.f�<b�ռ�:��u2r�x�❅ڿ��͢���nF	���A\'��$?�LnP%ˊ@D�WP˓B]7z8�;�pq)¦�0��`Y>�ps�������G�uO�Z%& ߽g����:��\A#~�)H��˅���p.�Z�t�9p�lW�B�O��	���|�%uZ�g�vt��V�U�T�ܶ� s^�_$���$���ߡ��s�3�&��K���+�:5�(;��~�/�D��L��Ϯ�T������0=�R�z�-T1���D�����|ee�xr.��r ����O�^��gHT���������h�W�����+���2�_g���@��K��t���9i�B��-T%�������{�{e��߾��6�#�~��]�ܱ�����7>Ž��d�7*Ɠ�}[�������Ys�]{�X6+q)?zZ�Qn��a��P���b*D�2��D'.Q%gkM1�����q�ABo~���R�X]B���|َ64�i��\z���A2B�z���i�@!!\��q���G��x}�:��{r�j�R��l�����g�%��u�H���$zw��>����^�R@c.dB���ح�D�9vV%2�9|{W#�r|{�wR������'��+���5B�Duob�͇0��Nk���-(g�|���6&�#sJ�b-�\]��r���G�0�~�	�k���(
�hp��G09�XaI�*��ȧ�-���)�|�@�s=q�lL~�x�����~�RU�! Ӕ��ID;�{������1�r�}�y^�p��ѝ&�,O�;�AM+����oBC��a���匾������Agj�{E��,�q2��!�t)��&��2�#� ��	���6�b�+���0Y��$☽�OEq�/r��uҸ�I�/�����i.ӻ)��іd;:J̤%S��M%���\Q@ȀaS����l�Z������.pS&W�3X����֐�[�h�Iq�isӚ3�0T�Q��UH$��T�qd^`
�(���S�};�Jb���AI	��W�i��ۋ1_��Vܜ�=z�M:�eU]LH[Ga��eP]A*�$\T���Mr��){�]&k�������;	��9S��C*����X�%�䱜|%�����!=D!ź��m�Dw�z� /�u>2TN�u[	uǸ�w�fC����N��NS�n�jG6��/�i�g���-�X���~�{#@���V����3
�a�9:��*�߁�r	�hd�a6a�fcv%��R�,���K���q�&�h��cĀ}y�U+\6��R��K �:�d�s���"=^�Y3�\����L��ʖ�4�
�Κ"����� ��/�r�7zե�w	��`�"�.sP��~+��Dx(���>�����P�|������y���M
6�R(V%e����IF�M6�5�}~;�� ޮ�j+<��m����a����O�o������$+o2�a�l�K�[�[_�R[[
���_ǐ��/#�}�����{�*��eױ��s�SK��ܜrBgyTg�z��)?S4�B9��Ę%�-�F�d�,�g""�-!�}��T�A=��d^��<9���
ӲR4g4��&7k�in�<�D���Ncv���ۏJj�e�.�`��Ҿ=��Nw�/`��:�J���S�5�W>���
���'eZW5'�7�D��ڨŅ��MH����z�ۂ@iz�C�cH:X~�"�����vQq��l��K�\���<��@��Xe+}`#��T���E���������!�B��C8���@� �@۽N�������+i����yH�E��t=�(�w��Z|��x��җ�R��E>V��(fy-к�q�>E̖ʚ��X�fA<C�2v�N��_)�W��Q�p��7�?ՀT4�dh��Le��v�Q�p�9�ˡ��d��6	��U|�u�'ZY�4H%��j��+�Œ�TB5VS����u/N��s�O�HݱQ]�N,�Ͻ�,Y)��bʢ���lRl��o:!s�/XhK&�;h�abM��Y��L�!`�J��*:k�{ل�P8W.��yp&?z�|����R���u[�7I �o_�k�N�6m~=�����x�&�ls���ՊvQ� �X��,��%3	V�&9��W���Jr`�J���Àp�ͫtg�����D���~��J�76$y|�ǜPc����K����v淳���}�L+C1���-���B����߬��;�ɂ����C�C=�|����#pL��3�y4�L疵�e=<�OGc�g�M>�`>8��Ex�L�[{LQ�N�.��	;�!�̉;Q��T@^�7U��O@`��1�0�D�0qP�㛲��h���]�0��ۺ�҂�Z��1>�O�C�hU�����L�K��?̹�+��h�6�⌟IoJ�M�����Hb@�N���<Ǘ zCTH�4�h��	��[��5��d�^{d0� �^�G�S/6p�SeV �U`�=2QUV�e�n;<I��ꚬX�@O�J�E��0��-i��l�{�}M�(}���LO	0x%%��gr�12�7*	��˞�^�Scԕ�w.���ǚ|Z\]j;C��D�Ǧ�X�8=��t�y�"U�D�C��Xt����l�KyQ��/:��7�֨}\K��~�������|K�[� �E:7���4 &)O�������e��\��F(:_��-�[ʭܱeX̡��ZQ�P�;ƱBw��K]r'�U&h
;,�G, ��ҵN	�٧ t?��ı�9t��N�xZ��4�8����p��P`�-�G�O�����R^O O>�R/��[�jl��]�Սm 8en�4��JUr2��l�H��aT�{�@_zX|:[z�>��
������~�
~���&փg�s�[[iA-�b�֤�Lw���ll�l�3��፹+�0�NN0�#LQ��}�!�e�%���h�������<7٥dp���~Y%*Q��Z	M����fP��O�1$��W����S�6��"�(!�۵Fa�ix��:����5�b4ܣ�eW#ȗ�M��Q�Vt�j��&�*��^l�Z+|�T��1�t�p�2��jg�ћ��wQW��a�����?��^DH����j&5n��0uk#3ªb	jєv�,�R���i�d���tM�Fl]8�y�u�V��<0�LL�Vj�tA�~S��v�g,�-e4�+cU(�.fF�ո�E��w�޹��ذ}Έ�c��̊�B�}��_:��]ԋ�
�p�����^Ӱ�ç�x�f�7�&?�7�'
2�?�.Uj���*�?O����q��<����_�O��u~�������^��f�U��+�d���US����!հ)%�1xfր�Z�Ͱ=�5��a��I����26)�N��S�BX(v�M"�Z#�0B׫mೀ�� p�٪#Ii�,x/1�]�D��Jh}5[���}5��Sl��^%:��lf�̤C�����f:�o^|�����;z��B�	�
�f֭7�nVv++g�ϠvG�l6(�aL騇`�~�k�Ğ�Dw��k2�}�3� ��خ	�z��7E���e�ib{�� ��W���(�M#ھ<���'	;yAƎ'����?�9�<��~H
z�	A}g��	Ȟ�M�Ad���7���E �|�����O.?�O-ʶ*��l����D�evg�m{�N7�kM�|D��i�ǯ�����\����y��m��(0���@�R�]�t�{W�F�A�c mh4'	���~c��!���N���u��8�n����$ �&�5hS���{*i��I�UlB���\?SŘ�+�vV�r�z2���"�G��[-I��e͸5:����?L�.Ȩ�����h/=>��kF�4�6��P�:{�_(��~R�!%y����?�;B��6�NSe��a:�4PT^�[x_�
�Ɵ���q��.�3c���U�Ĕl���U"�8z\K|[����=�� �G6eR�x�؛9/�q���
ѳR0�cL^�:���3Q��l�>,O�l��QAm��!
I��"5�J��X <���K�W4���Hi���?t6;��~C���_�[*%%(X	0�{��_��!!���&���֗��cs��f.7W���ubD������;�
��`�K�8Χ��U�����><�9�D�D�M��t3]2���V��'�Gw���AG���(a۝u��ƕA��f`�"�^��仠��9�x\:���v�ڹ��y�S��}Qɤ�������\�?9�M_��7*��5;��(���Qq	�;N*���~*y"Y�%�Ÿ���	��O?��|��u�����s�M��g�e �W{|�X��P�f?PKZ+ϔ-^�+�I�wA׆�"��9�B|��&m;.��F���T�K��JV?Q�cR؜G�.vLe �T��l��܁��E
��Nބ�%��.���;I�����SG��`�v/1��
``��kE0�lf׀g ��#��4ױ��lԞ���bWu_h{�J�#��"+wA��O�n�� �%�=�~e���z���A+��u���itv��M!��vP�G`x}�G�#DZj�BR�@�LhD``)�k�Zi�O��_ʂ��!����2��&;$�W���`sG?n��)�CB��{�(���jj�V����R)�+`Duc�PZo� ��#��x��s$���~��!��ql�%��:|ɺ��lmڒ7�C����y�Q"'�T�S���bm�ҩ�5�f���R���:����H��Ó�R��zF�6a��_bM���U���|�m�1�"ᰠ����5)*
�)7�p��������à��ʧV�N �� �&X�� �B��#λ�Ø7�~�nM�ɣ�#�Z��e���'�rs�	�\�c?T6�O���C	�gͧx������#.��C�f�7Z�N,�����NGz�'X������p|˲D����9_'��'NhSJ8��
3��}�w�w�M+3�s��-VORݔ \����-|#PeP��!&\DI��\[�01�0Xa{b�9�yt�%������s�Z���hr����ޓ�X�EX��jE�<����/k�:+�Vy�d%#��|q���"<&s�x�\�g�)��X�1��u�S0c���C}���@(mY�o�.�{34f��lJ�v�+��R�	����NM�l���	-����cD��֘�sK�!Q��~طlNͽ�)D��Qer�F��Hlb�?�S���%�v���?�t�~�E�_������Wc���A.�$�
w�{��W* �7Cߤ����r��X��ow�J�GQƿܬj�L0ߛ`*�i��&�I�&�_��{����c��'_���g����q�/T���P,X���H;�75 o��W�9Q��q� �UFm��,��g���a�ˇ�/���[؃��2��u��Oȅ}4���x�n��녓[���$9�Nj��:'���P3O���G)��t����~L�jy�w�`��;��@ʓ
s$%�T��M��i*�=~��Y�V��x�~qȉ�t�o�����@B/�m�ӽ��i�λ�V��k����W6�a�>/�O������+'�TX�hm�������ρj�߬�	v��'���S�U
ʤ���\��9Z���^{=|��Qĥ8gB�/ғw� 2�Lj�F��&RY�(G<.8fxd�%"%/7�oD=��	DX���W�������{pt1Q��{[�t[w�K��==���݋4s<��_��F�a@�
��,ap��kAL��3Z�}�ꃑ��Rh�C�Q�2�O����=.���ǂ���Oo%.[4�D.����e��M�+���8��&N���Z�=��Ӯm�_�*�ޑԢ��5ܜWL��E�n:�j�tT�2�(�I�d���{�88 jH��!H8�z�I㋽p�7ٸ��Z�ċ���T1)���u�t�NXr�+
�G1�}�$�<9�3���[���[���*�34��Yȩ��k���-�hj"�g��>�8�L��!%!��}K��`@#&j$����-2>؊A�F=b�C2>��z_a�S���R��LR����f��Oq'�n�ɤ�6�?�^
��z��=7�����b�+Qhp�r��Y* #'�w*#Ae�9�6�.ĉ��[	�� F��A��z�$nX�[�L|wN�ǰ�����1C��֦�����I�4�R��;�EW����9Qh*M��[�|;��n�����P��a���Ur��Ol�~$�)w�tC8�v~fg�8��b�ɊUrݢg��NiYk@�8�� �S�E�(�z�(ѭ'/H��TǤ�80�0_6��~���̽���g�+��Xo�ry u�E�b�W����$r"D���o8z�!���r����� ��}FĎ��\�]­�k�@���|B�(ob>�\���.
��ГS��	s/���T
���chR��iO�A�"�-�Ƶ�_�ѭޗ.���g7wR�����{tl�{\Z�{@�����;�s{���hJ�����W��q����{b��~X�*�tC���sg�H�+z�I�̏�� ���/�o�Y�O�%�j/-m��������5}�ym���V��:5A�5W���3�`iµ����>��P�#��q2A�~(�Z�N�F���͏�����^}�D �&�� Du'1Շ7�0g�Wn���s�m�������\�7G����Y�PJ�_ـ�~�a2�W���������3*�{v�=�#���ϟy���ā��~��C�C�_���Bi_ .��Ts?������p�F�J�����#w ��Y�/qN��I���,^���" �5|4M�4欍&��%�w����hT�;�B螷G��d��u.�����-T�X�Um1h�~��6�Z����J���@���A
�6�	� 6]�͹���]��k���(^��(&��t�}�hN�w��1�[7V��?�P@
�Y��u����zP�Z(�v�����.#G����C�>a�98`������V^#��Zx�{XބX� �fX	����K�-l��kawӵ�9�I�q�Vf�����)�;�Tx��2�ۛ��[���*�I�p-jX����2	�?�-h��̥�x��JÇgd��O�H�%�_Q�@�C�HR��'�H1!��h�������OC�x�����0�JyȆɽ�>`9���XYJ@�Ȟ��6���(�UU����6Q���5l{��:T�����I�������J�t�+2�qY�x�A���9��k��g{�� �yV`����g�I�d�!N�4�K6􏗲���
9�u�<���o@S���
�Y�_��&�iQ/ 9��aQ;w��tۣ*wƺ ��NIM�Π�ç��N���a��]A�kpF��?�r����6�!�̌Z8����E�l�'�G�ΕP�`7Q\�(��ęYWJ#�TH;�Ti��ؑ���e!"��:��S$��e�zvxT��;�}���\Ȁ����n�~nf6{�j�����6O�$<G�{$���͈7�8v '��痨m^�wk��p��2<�/?L6����Bx����C?a�*d\Q��V�E���2���-/K���iggLm�%b�_ ׹5O�ngP�e�$�Q��o�7zwp��,)��B�.(��\��F����v�͂sS?��:����y:��Z���R���]���-����􇡭aᘳoC��M�Y<�^�t���/UðF���8{��@#N����P�|���c[�L�Y��j�n�����w�[��y05�F3)��e�v�NX]�t�JC�Sdri�zZ�)�eQ�\|��B�	��'%q_[6ձJ���O,�Bi=�;j�-#�AO�f3��z^��7���cUBr|^6�_s�V+�X���aH��c��NIyW��1hY��q3�f�~uțy�g����쎞�ffGp�8���u�	������;p�gY2MP㸶:����Y����J�i��P���� �c
S}��-��Oyn�1���9�*���?Y�~��K��Q�p���R0{�B����&���`W�q<6#T�a�Ι,K%;:�M$PO*n>��i1�zi�o��Nq*T&�
C��Ԍd���>�BF��D��u?���?9�L�F\���,�1.Y��W�h�K0Y���ʝ�@W$ϾX�;@���"C�"8�v�NV!�f�O.�\7��X�y�H�:!q��|�5v���o��a�w�o�/:9�zy��Y$�F�)����ݛE��e����І�j���R���9�� @Y%���F��4��=B!�H�e8�f�rqT�oeq뼸'���9\��v{w���=�rʼT�z٪�̹
�I�})\���P
;d��{��A��\ޤ`��Y����,2����7e,2Mx����<L�r�]x(nk�Y7�K9K���)i���;����{����c|ׇp��^'���pӖ���X������ÞN<I�U���Dx���_L���m"BI&����|���b�C�b�x*T���!���{d��ka���Q���/�#2`��*d���w�P�(%���.�Ig�7U����I�~�t��\�P��h���ߔ��s��p&��9v����YV�ڝr��z?���ō����Ʃ�:ep�����Qș�!V=��l�ءb�dd˂��&Ӹ뺷��iA@l�Mr��;-��f6�K4�ڑl��釚gL��`�LҺ��DJ�ٻrľ"�f�p�2��q��*>��
0Ĵ4��9Wgy��)�`��"0��i}�<�b����>�*�^���>�MῡM!����
=A`�;��E�3�Q���Û. ���8�8f��j��S&��H99��b�@]�˨a^^��~ ��6g<9w�����ũ���a4*�<_�������h~�\V%�~�'�D�F}�!IRg@�D� Sfc����x8o�(?�2�Z����1sW4�����7N-�섀�78�����` ��1p��.7��5j�hh
�W#�(y���c�
2�}�c5Aʗ��^�M���"I�Pg�$4;��$�1:�*�r��;�jR��H�$�Ty����Ė< ������E��t�����1�۳����aU�#$r��9�T��?��ؚ��X��ja�U��"�t�3�8��a)VP��F��A��(<��$���?� �T8��48#ec���aAd�d��]S��s�?#ˤ����;~A"29�/'M��R��.Sز��������!7�E�*˙���B�E�ͮC2��"ڦ����K���z]-����C�uF-���©f�E��]J��!�L7�p[��/��L�6=��'̠0��
]8�x@طe��l�h�"��B3��?M��Q�"�ԧ���!8݀$�V���^\vb��r��$��I�~3v%s��,�v)U���{>7C�Y��:�¸`^��'��|Ӧ��o���2��W�2�;�q�w����@sّ����Ǟ�E����({|d�%�h}�����+�dm��L0�}�FP��X;�JGB�k�0K�j0��P�N���YWF� l�]�A��|�Q��.tt�,��N�G��-�GT'�Ŕк̶v9^�� l��]�Y����9��?���E��[kz; ��&��7�'�'ⴔ��/�[Wq�C���� �0Ҽ���[ �i�Kk}����NL��7x-���n`I��I����B��\F^��+�&vUD��+���,I���s����Q���4�l�� C�Ƣ��:ݟ�@�i�m1{���P�,3A֔�ڂ��p3�b�$���.�a�-�(#�)ҭ�Kf����@O��y�oT!��ʘ|���|D̜8�` �Wa (�ښ�R�ڜ��0ɷ#�U��L�z*1;���j��_B�<�G�6��3sC��(^e�����s���K5��`Bܢ��@���v�_Q�):�����������sO��8�'�f(���,ʽEЮD���[����%� {U�W������2H ������� %�?�
^�O�Fl��G!�Mݤí@�D$diC5���Of��su_0Xc�� 顮�ϯ~��G�CQ&p��&R�X��@�>B�y���i��&,+�����'�>$��S5ӑwP�T�����e�P�Q���#���kа���Ȭb���e!W�Hd%��raÅm�����%൸��`�a��{]��5�B�T:{�ђ�B��|�돠XL��`nr��L���� 5"�Hܣ�	��j�/㛜��b�:�����ˠAA�f��򫣾����8�e'�U�N{$��xa�����ه@-�..Y�Ͽz�[�j�6ʹ�m&��J����)�~J��?;5��'/��~���(L����Ʃ�i*�ff��S}�í��ݘq�̼��	 �r��<+���
��\�L��@-2{���SNt��1O=���((��sٍ�U@`�잯W�e�,�I�c8%��9���jho���؍����Sc�8..�樃d$��(yX .!VOMɸj��0��.c��F@��� J�Gi9�%�Dm<�V�F�Zg|�6�ٓ�>�ЯT=i�x9FL�/B��r>���h��7~9�,ݎ�$Jbo��FY��v��5q�Km}~�pe�84BC�4T�b��d0��X��ԙ$�4�Q E�2
��w9o�p���x��]�35Pw~{dˑ�)+M�o��'�u�(I�K徹b��g��*丙�Ha�� Ǖ쮐���5+?$k0%H_���)���R�λ��4�ޒ��]<�ʍ��Ռ�ˁ�����Ƙg\q�x���e5�3�D�No�%@�B�Opo|U��ʺ�΅�$��Ġ�͛d�j�o��oC�4��^��>`?�^r���.6�8�-&����M������dv�F�-~�3f�Ѽ��*�r�Z�́���C��~��ʼ�Wo]z��E��5�z��ݿ�$�ƚ~cg͗6�9/�&������B���~P��S�w�fc���XLd�x{�����ʇ�k���ւ�E8�Q��fx9��R�(0�I�#���:ˠdxLYlz�j$���uA	2�M�����¡�]@�=�*����o��n���X�
����|d��|�a��i� ��2W=��E㥶��8Ý��$d�W�>̀F�Bҁ9�GʃiJ����	�:3�	�f�G"��2�������4MW�G(�C�V��x��Sx�S=�tfȨUG�H����S3�1����T�,�ԵDB0q:����K�Bm�L$)�s� R��9�����g���?��1B����0�o�w�ťV]��f��c�$�(����K����3 70��x��)O��>�ہ�7�Y�n�,������ )�E�de��0wj?!^��e��ȩ�z4�O�%`>���Db�{��$�:Ͽ�*D���\ݣ�i�mx��w��Nזd�j��9�1 BU=��%|����X춄t]h��y����Mj[O��^X�_�M��W��/�LlY��hUf�ɷ��|.e�I`�a�Z3
,Q�%� �#��)���8s�E�L�\Ô�n��z+h��Gj�YO!�������^�	�����j��7�3�98Po`������� >85q�_����pO[���r�5O��9	_擒��W�,qK6�Q�- ��ئ
f8��;�yH���z���@��0���	j�_�E���g�����d�l�Yg�8�_�"����W�v Ui�N�;�֐S�k2{�[ӏ05a��e�g��-]��{EEH�/zp���|�C�o-3�ߦS�r�.��%r��Z����EA���s��J�3^MNt��n��e�A�S����
U1'w�a}�4�j�Ŀt�i���إj��"D�CH�_L�0;���И�|�ґ,:8��@A��.��T_�;��M��9���8Dm���7�w�(4��F�LX^��qJj\ޥ�_�*�jJ��|���U������ ˵�v,�h6��"W؛���Gw1����wc��@rNb�NN�P�S����G8Nc�-��?��?��U����L{�>��;��#ju�Ʀ�h��+�9L;����l��̸�2��7�s���H8�۝� U�]��>$�ls_X��Z�����eH�-��������wЛ�d ��L$-}�����Y��p
�ҽ*kB���������C��W4�ޑ�ɖU�C��B_���6��ϧ���he��oߙ^?��W�RvŻ����GAPҟ5��~n�JI{1L�� ƚ{;!���M��e8
Q޴�d4�XR\�4ȡ/�n� y��}Q�{�	��Rɺ�9q��y>�p�0�iE�I�Y��,�3�T�:������ڡ'�io��3�9R��Pл�jݟ���7��F��|2W��<}�m�)�޴���Hȉ;��?Y���&2�z�����сo�ˈb/c%���ڈF�����bߦ.	���p��6$�{5�*9w��.Hoqh��l	��緦%�<�b��-�#ᙹh��Ln���մ�xv���z <�\�������-΢"�8���q8��[W0)r�i�s@������1
sD��M)�����w��E]�$+쯻cc�7^��?+����r���l 3UiͿƩ��ʙ�-�a����Y1��P:�$�A��N���k��r�fgܾj�Gh
����cԈi�����c��Xƙ����r:�ۆ��^&n���af��8[B;�'�@P�d���~Йʼt���~1	m��Byf�n٬Ƌ�Q(�8V����]��}o k�l���4[�!c����b�XRR1mn��U���,C��K#�Eh�7��~���]��ߝz�i������]:��j0�˴ju��Y�u�4rw/]AK�X�\���z��J�u �Z��D���j �o��,��/ǈ��ʮ�H�m-���ߴ��]Q�?�Uᶜ}�x�dn2g�ۼ�a_�,2آ/~|�#NHw���p��kч6�u�r��M��`V ��'e��%{7�6��C�-.a.�޽7c�X��2�J��1���>ѯJ��N��SS�n�{�<�o��ܒ��,TF =�El:[8����M�$�1�e a����<��Dk�g��n
���y��J,o��h��|}����������<ho#d@���O��Lv� J��������b�;�b
��g��l��W��Y�Kq	�	�a���)F��?	��s�ũ��IL3���gS�M�� �� �8���?�a�k=Q��*B\��{i���xu�yL�x-l��S9�)�j�o��	ڟ\@�>9#��>Y;��;-x�D�7�������s�{�؆g�d���c�\�;�\I��C1T��(�\����&!
���isEe�����48��:���-t����O�ɡ9J�Q�+ �vw�-;�9�^�h�
�"��`�)
Do�x��NX�p��S���h�^��2�*ƈ?8o`��dV&�S1nێv�g��'�+>�����Q�Iˮ���]\��[y��־�m��"P���9x�*Ρ�W3���e�6p�+ʙ�������Q֎x�J|*T׵f`�D��XGz}}+*sA�6�ҏ\o���\-vh̏�}օ����})����,i�d�(�0�O�}||�g�i>�9��Rk�q?蹔l��#�����"�ŧ�)���8�]AbH"KT��x�eD]���;gn�ҧX�c��,L�pQ�$�˅V[��k�5���&5R��ֹ�`�:�j$V8o��Ҿ�9>���v�(0���H>ޔ͵,+��U�U�{����]ײܟ��G���{���`
�xv�*�S�ű~,,���z0q�礧�f��}�<�]����ơn�*���`B�Z���mMBH�#r��>_� �0G�|��-6�K�E���(��*x�,M塓�"E
-	2C����u�>�$~� y��ᘴQ^��9%��*��ͤ�*�B��m�}���ٷ��Uώ��^s@����Y�[�Ex-)�Yoy-lJ��;+sv�����
n��ף��
�$��i��)�!��L��h-�=\j8U&Α}�#Zx�
�v�DU@��򉍃KI�o�CS�&v�099��@I��GH.����'.�]N p��T���n�J���hS%T����t��� �_���.�^Ί:n<����f����VQ�5�-Qdj�P���1���T��}�����Y�SG!�Z/�;.��ăPצ��
y�Qp���v6��dC�d͔$�2�Y��[����x+������H�0�в��ɏN��0�O[�L�q�M��B��Pԯ"Q��g5?:�X&6x���q�U^y4�JQ�}���/ȵ18밢(M��t���Q��6ݗt�����OҞ֪2]v~�Š�k�e
\��.�2Í �
��A04ʮ����51�^���h����/Ƶ���o���g�u9W@�)������6�W<�1"U��OAJ�s��U�W�˗9�۲�q���E��N�Ĭ��8�Ydqp��_T�9�����s榫�D�@b��®��#����\䈷XnH��v[4lf(���>"p�J(B�l�O��X�®���׿V��᪉y��(`�2\wZ����O�u����h�-i_�KZ���1+ط�vǯ�V��=F�1]M͛w��޸��wX/f�\K~�ymQ./h�G��n��Tlsr	s�>G_��H ���*�����k�g�z�"/��x�Ҍ�'��|����ڢ�ѹᖛ_��w����T`Ie1�2�É�N�@jt0c�	�d�9C�g��9�ܘ��[d2]���}���67'���c��Td�ƄC���]Μp����ahJ���E�[/(o��?�=�j��Aս��X7NvNo��B+�W5rS�W�	q�&�{�����bNyA(ش�4�pƢ����7�`5�)�=���j�;�"��Zڔg�?Qp��;��� mj#¦���3r1�l^v�uMo�Ճ�U�Gq�QEC�6$v����k^R-<�g&�=,8پ�Z,���$gLnD�RM!�ۄO��r�]f�z�j;�	�\ U�~�)��8#����a,�d[�An��I�+��'ϠJ��Y�������LQ�q/j^$%����+PYL�.�-6
Nv0�"O��G\C��d�==u{����yaOV:Mӯrҗ��<��}�U0�э�K�N�fD��wQ�q֜ꛆh����mN��]�U�`�8�T��*�i$ ���W�+OP�j���c�ZU����i�Oj�;��}BD��ԯ���E�%	n���t3�(B�Jb��2:�
O+�g���	z�n� 4̓�����2N�����%<��������S��|�NI�����"(寮�m��]͑�Y܀ ��d�ȟ8Ǟ��x#�x�Zϩo;�A�V@�n�m�:=�kt���a�. u���av�T�Q��8};ւ6Ym$G]�B��e��1w8#�d��d��?��y����oJ�]��ݞ��i��XV�u��97-Z��s8�h-��'y1R��ks1vC|/K,�Q�(�G]=� $�Hu���:�wC�M"y$��",F,f�"�'D,j�ML�zd�BFm��*��[6����v�`��$t_2�٩�r����� ��,`�T�2���)�BS��e��6�5p�	�$,�|wa�N�<��L�=�C�~z2''��:��b��Z���DC���)�J�p�����ħC�C6�Ve3���UdO�d	U�A0jj�'pdO#�:� �����m����:���Ă��W�Ƙw�Wn�C�~��>��Qn��
{����
�`���aE��	J?Z��{qbx�Q��9@uQ�:jI�ؗ�>��6�/e�\�R�\���{�q����q����W�%Q�`�J!B���Q�J���pj�v�P�����N�oE�]0v7�_�ɾ^7��e_���[&|�������^��b�l^�XaS
�\��֤�g�C�o�9βv�:/���p�b�p��f4�L�m�ml��7�ԛUF��j(��A��D?x7�w�C�%� p{���1W�T���yQ�������>�z�B=V��L+*�N�Di^�)���m&,���2T�o���Z�_���Ɩ��]-"����Q����Z>���[LCB�bX�7=���M��Ϊ��)ƀAl zN|v�(5/���±��y((�L��������JiH3�XN��wSR��Y�a١d|�F�aj�Uٯ8�VZ9��8d�s�~��r��n-��'�7b��o���Ф3sC_*�؄�U��]��;�˻/�h�&P��!�'(J}"�gt�CI1?�Mf� ���1��V=�,��	�@�1�*C�6l�Gl<����A9�d~���`<���v{SN=k�w}���<6��I�Cs-���/�����Mk�P�s�Z�����5���E�:�P�x�ơ؍G�����#��VLq�� ��s��E���������ZN\ԵUѡ����L��G���%���
�b�'�U��1x�P����|?p���tO!��
I��%�8f�ϪymȌ�����C�|#@�쉰4�▴�~�%`|��.l�64U��W����D޼�;AsUW/�_ߘ�8�&��~�Y���3����I���0�^>��n�+�|@0�*h� �\�z	����<��i*��1QB�r���,d�a��;�d肛��T�w]�K�`k[X��
��f��mȮ�h�;w�)dX���z��������o�ռ�wJ�&4e�k|�}i<�kd]����H�ke�!&y�VQS�am���lz��H�r��^pC����y�W!�{�{N���a�������rs.�mW��i�g�&1G�wzI�#0S �L��3)Hܡ�4�k�O�j�j�o�^�o M�����| ߋi������D���eS��z��Dׯ�d��UF &��(A��y��H�����0��%��?�&�kQ�g�^Z9�B�`xV�M�������� �z�//'�a��P���+:s��:h�u�� q�S���$]��F��B��^�T���\�H<o�`�GT
���N��j_}q���6v;�Q��UB%�\ܕ��m�z�	�!5�kY��D�e��(�Q1���^�:%ۢ�
�~n,�KQ�T�Zc�ы�^��nmD����w��HE����ғ������&���z�� �7#g#��*+��)a��y��Os1�Cvs]q�����?��p0�ݸ�X��v��B�����K@�!f��9����﯊�He?.#qCUDЉލ����g�4�em�����o}ΰ'�r;��56�W">�e����em�Y`л�EΘ��2'!i��Z!����׍��? J�e|�I���@���0�<ԑ�ɰ�JTX��w<���b��P�)&�F�*Y�NkP	S�d�F���}��-@Kn����M��we�C�T���&�6讠�qN5��`ZB��W�ȒCyL#0O�&f5J��1Kr-�~6�j��#� ���.��ǧJEsm�O��T%�M��|o��^j�#�I�M�5��Y5�QG�� T-����,�0�'q�V'�s?B�IZ��d�+ؗ�L҇�A�y���%��:�J�a���v-٥y-$�d���~*�!�|�i�+��[���vE:+|����٣E��-��x�_;lӞ.�%b����V���@���sv�������хq���׿=�]8M�0�J��J�C�&�)H6����Ke�߇�z�R��
�w���[��O�����I���䀱�SI�N���"J���/ڑ�<ݵS}ƶ�@A�4�[1`��9:~�Hxw�\�I�����i=;����g����J�a���vI� FgKc�����o�P�b�ݖW���ǉ��a��[�j�~J�:�b伝�A�u�L�<�3���0
��ׁl" 	ΟL���˼W辱)�5�ܗ��x�S�7�e҃�X���v1�Й�)C�m$�.�>Tn����l�q��JxlZ4qǢ�hC��#_�����0wU��"�]�v�u++����Pu�K@��dFT)��I,>m`[��H���? +���ެ���O~���L:7N�����0T�-D���������~=�c�a�P�.��zCc��2�2F���;o1RY~�|�/!����\�hQ�|���&8�;D-d�dL�kD�:�����X�������˶�~}��N��D�_dk<�*9�8��㚋����4��EB4�`&������;X0ND��8}H�*؃�W=r{���~�"E���]�������Y��F5�2�w܋Sۣ=�����r> _�v���`�'�x*Կma��K���	�v2��90T�$T�)�U��msy��WŲp��պ2X�e���|��B�|M�)�Z��"��yUp�҈Q��������I�o�G�*{2�^j��0%�v���.�z̕S��sh՗���]m�L��k]M�e>�>n�;8���Nɞ�4�s����2�:�~�(]mƞ"��D1�
d՟b�0�f@��!n����nE�{�0�����T)��̳I�<��Y����Hp׷�)���&f��ǲ���rиz^|��qU�Xܺ�)M
��C\K)|6�<X
D#��k2�ñy�A�yh�:.�V�T��0�U$�6��{�瞴������1�g]) �]��9�\+~�^K��,c��`����P�tIo��P��TD�*h�<�N��X�L��_���6�(�Ud�x�s�M�:km���-��/��M�K����fV��T-��q�~~f��U�l����%�a"�yrZ'v��F� I�G��d�3���p;�Ty�� ��8��y~�f:���RL&|=�Qw?T�x���E�6t�ٽ�����K���H^\z���H��s�a*r����Xl�y�ޫ��B
����@3�b���T�	'�Z�����,�E5�w�չ3�i���/��u��?2dB���D�����>�K���]�٩�IG�7�aAw�K���������~�..OƢ�m�#�ތ��WKGL����칒�($K-��V�+���	i�P�x�����ӫ椀E�šN��{���Χv(�x
�))���}����P�ʡ��w<���YD�l��_�3|�����+XT�nkXf��MwR��8B*�d�:�flTl�Q��)#�bt��
��#"<�/�DP���߾�3���*]?�fL�3p��7�ތ�̓=�A=�Yy��Dv���!4Iu���Y]�������n%��g����h�g�d.�G�ub_S}ۓ쪿�2�VJk���j5Y@F����"}�h���f�{�mЎ�i��^6W�^'��3��NB|ƩI���F����`w|�6f�����v������|mP�G���*;
�ܦG���].��8���oa]Rȓ#T�W��:؀0cK0-n�>I�%�>>�Q1 V��w����b^L������a���{�¢���G	�`�s��`1g�������*!�Ǻ��	�a��}o��e�*��Wj���䤗�^��>P7{���\5������.-��#��K���j��uq.��|�E�C���Ce�BH9�P�вS�tq�f|!�s��#�Z���ߘ��&c���# 0�����:��T�aX��Z�*�T�M?c���D��h�G�O���?cr�ԫ�l�ЋJ�H�=�"4n�[�6�#�P�~ؾK�}�o��7I�W�����Bb6�ݹ�7���i�9|'v(@��cV�C�֪�O�y�4��͐?b�h޿o0T7z�  xHt�[�Х��u��3|k#�-�y-s���v�@�_�Ll.iJVb)�:�M0J���y�EY9�U�j3�8o/M�s�.�z��m��8�Ȝ�O �D[�g��"�h�|��FE�?i����Y��}?��1c�ȏa��C����^�]8��&�u4y"�-�^`���������������u!�^6�7[��OV��f�-D��:�_�s�nCv�l�6�u �D�c7�*W���v�;���CbZ9��{�1l�0Q$־�̪�歑^g��r�� tx�#����|;#~HU�)�Ј�a>�
���R���\�f�Gj�V?ҋ�SO-����������#��!v<s���j�9�K����r��'K�������e��3�s�h��(�q2�ʚr�a1"e��@Y�=F��I��.�TyP�e�1.P]c�AB�1Ր��9�N����;9Υ��P�vU{��%Ȯj�N��<N��#�5��5�0��}���u�AS�0���Q�M�-��7��P��'_:������-���T�AG�҆�A7�?o*�v������.eFZ��&�*ފ*���q������K����8�Q����=�K��P���b�A����;C�8���̉�n�����2���[��s�K���
��p3�e/�A�����~�7��k�1d����:�� $�Ͼ�Թ��w��K��%n��ۛW�╄3�%R�"�ѿ�E�r�8U{��A*�%W������iKj���`t���R[�~�����IOp�qT�V�#k>J�#K6�Y��Z����a@,��ZE�5�3 #�ӛ���)�5�����ҞP�H�g_��E"b�}���$���[.bǥ��=C��6�\~j�4r��ҙ�f&=���\t�JA�y0TZ4` �t��m��F,Qg��Ag�]$�[��D��O��n����P%CB���K��^&�9{A� �{��2n�#o-�$}^�%��+�#ļЏb!���%����.��|ɨ�M��h���0�d�)�	j6O�M^�Ԝ[%K��m�r[���T��ޓ��=�E7j��x�s�R{���4q�(�ZO�z�Q�Zb��ţkd�4@ֆp�x|�*@�d|ȩ��#�sC�Z( ��}�Sz����<���Ȫ�Ϊ�C�t<&�;y#\�YŰ)�<�h�����������_?n ���Q�-�|ً��յ��]��+s�N��ofp�=|_Y:͞����ԯ��eZ���g:i/�m�8U&N_v@!�\������@¦v��렋,�^��Kk�@
�K�rV�����Y�41�WS�L,N/�-��1B��&�B��젅�xiT��A�˘�,��F%0��䤨���Y����Ag���(��?#E}O��p���wn��D�:s�^8�M���"R��#��ռ���K�ߣ����*�.��L3����-��l�-!VԞ��<�L0Q{�ۿ��~�b@��g�ꖫ�F��}�Ġ1;n�;<��E�2
	j�z�N�@��v6f%�U�g���t%�Uzʰ�"��L﹕���Lė�˟&�?�T�d,��n2�:T|)�ncE�a�k��g�Y���"�_,�Wb�1��i��'��%!3'�5.�T�ۋ'B�1�Y9���a�x'
nۋ���F�X�
�^�l�����z�6sǘ�F�a�~��I�QT��Q�'Ͷdn��D�����6d����j[j���Ϋ�<�R��7�ίwT��H��k�C9����SJ6��5�e��7y>��EZ�H��Ê���Q�#���2�E�����K�;�k�-����¥�
$b9��`�8��d�+o`��!����q$	�<�� ����L$d���
������_bz�f�� Qq*�NO�}���Zf�$����=�����ڤ�������}��/$�z�ϚG����Z�cՆ6����ld�%��C�����H��k�{G^J�n��)@�d��+�4~�� -�hOBOf3��Z0r��[���Xj���"��M$<������#'C�f�����e�>l!g��@v��j���S�z�ī�
pwWg\��#S�>��g��?cXy,�e83y%ދ�ޞ����W���B�u�k�<X$�4�ڈ@O.��ZQ�L���N��]����� b� ���sw{�~>Fn"�O��)x�C����Q>Jh���Si}(�0:"M	���ฟ��$����G=�������TK�j��)����xr��.��������79��q[�l����V��ی�����2��
��޻�ӸS>t�y�G���b���h!�&m�Q�I_)�Pzx���7��̒+Nq����QG~��QA�?�p��U%N&�2a\�Y�\������+���38,����s�5��L�����cc/K�Ҝ
�=NÖ�����1g�q8� �l�s�iW[�E'%����e��%�!�eL�4��
�V�wM[��*̬ڈ�^��� ��/�ѢvABx��_!�"��l��~k�X�kaV7d�������"r���Z��<�	��?�A��C�0[��[����P3���m�������ϒ�A���ߏ�w"���ギ�eOE�h�	UR̰~���sq) Z��:��t�e ��Ϙ29�P�O����<�D�X�O��Iq��s3��b^��Tdv �l�b�j#ܰ�(n�����=����%q
x?"ZxSV�9����olT�oA���[zJ���������Qq8�H��t��ؖ$-z^��6�/	�B͠RhD��&Q��# ��vie��e�m��W�=O��h��!3%z��`*��1�_�����pȭ�g �e5̹ޑ�8� Lg�I�PA�A�jֲ����n��ƪN@E�4Ug1B��O��e]��}�u��f���OG�hl��Ƿ�;�3|��t"x]�FLΣ[4o��n�K�>���� rzr��Ɵ����6�3I��f�� }<�%|x�f� ���ːf�'wF��X��(j�2��{B��O�t�*"s�"�.�(8Jú�5΁}��(����zR��a�앹d����ܫ�4��	�Mo����g�<���U�?�D1��o��ke��tD��n���_���8��H� zL��> Z���`�9�]'}���ë�}P�S7EՀ��[=��=���b����"�9�މ�l��#�6&2�K��ޗ5#R8��	LB�Rs�d
��#��τC�]ܽ�/�a�8�<GmGw�[v�vv�LK���hK�W��ꠂ�1��ڏ��װmixLͅݕ�E��#s?���!�r���'�u�P V�wάk��Ywmu��&I8Y��^&ި&d����6�p7u#��	[�ǙN0	���7/�[Q��²��W�p�(�zG�����
p���|���%yP����,w��H�,��",b^C�T��n��2�l�1s�P���xS�o��\�~�O��q%���m��B=��/�V�l�-)ԡ��LB��Xbk���,�s�1��/%���'ϭ"�<.�
�<%|!S�$���1q�YFb��7�[F1��R�����^��c��8N.�Jnk���|8�~��m�/�o�����$x(,��03��Wd�����֪��v;����h�\/�X_���M��6ۛ�0Z^>N߽��݋�� ���3Jq+3��#�j�҇�5H~�9̤A2�m�G���sh��L�de����Y��rP����׷&&'l3��X��B���niUpy����a�s�!��D �$SYx���	( C��=����*(�BlE?�|��HŚ���ƪG�Q+�xS
5���C�o��7v�l~̚Kf�1�Bb0?@� K��48}�W��`����N�X�?��>bNڊ�G3�>_�-�)K\�_i%\�`lD�u.�o�_����Ǝ��N���_�ݾx�ݨ��V�Կ�]�,���+=�U�=1_���t�oq8��"�2j�QY�Ø�X���m�� <:���	#$0hY��-��k��OI�j��{1	ͱ�̫c-rS������)3Ƀ~�~���q+F
K�(@��R�2��oA#Q�9k�I������ch�8_]-o�I��2�Zh�z�l��U����DCA��Re߀���:2
�hja�����)��p��|��/�ܲ�H�d\[�LJD��1(%��sk,md�`X�U��% ��J��I���E����ɔ���
�����mt��W��2���@��b�