��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ�;+G;�2�̋�
F)a �*�Q-�٘9;���ʮrI�h�=� �0[����& i�6�Ř/�˼�����C�%�dR���m���O��G���=�����U��y4׀�J�x��~�tW�l�&Wj����Qt�Q�#k���y"0��ȼ�$����K��hc,�W��S�_��֎���s�D�o�z�>4<�0��}����l
Z���6��Q����c�[��a#aU{�a�O���Lf�p���G?Yd���?o��<��[O5�E��� ;4�`�� �`�F�4�#����!����˫W(ߚ݁��5!�4$���H�L���wM�.=�.̵���)��
	��� �'�TPF��X G����q^\�s�*�*�ôو��s(�6d�Ǵ$�#b��TZ�Y�(6b�Э�t ���'-�B�&Yͤ�d*�G�l����/'���o�e5�_�޽/�a����l�3>����7��>�ҙg*T_�>QH�} x�P������9U�Z:Z��tyZ���(�
�1>���O�a���[�T�C�cx���_u5nT�6�����V; HN"�����^&�ܭ���xQ͔9d�Y$m�_|lV�Յ!�ȣ}:3E�U<�ػSbK��ӷ�Ԣ���B� ǖ��(9���"=g����m�4�M9%]�>@1������;�}>��tS��c�%�KQ�Bm�\0'yb��Ч��{w�NgT�J} ���!��E�js��ĴX�ϫgZ�)+gvc؎�-"R~L��ߞ>B��a�>� ��馣Lv#7JU?���_o.Ҫiyb6K�Őj�kc`�}��u�3h�q��?
e|�G�JEx��`J&�NZ�c�$�B_L����u���w��'��������}�`��/N�#=O^�׸�s��h^�֤����C��Q�'���}>z�Q�ߌAL���2����lx��T��Os�����"۝�����IC���&����v�?a�7h9��LR�8/��㚷���q)L�8֣��^�ȸv���Z�f߄P�R&2ƈ$��	g^`�.'���!�<a.	2�a�vw|��:����T��V!� ҫ�!7h��.e��Υ��K6�����~��,�μ
{l��x,�T��|�Þ�C��A��3���J��Z����h����f�G��ĳEImr��ƨ�������Be��]ޅ�(�r�eI&yQ��� �XV�T��KQ�Y�.,��z��N˒u��*�?�aW��pʑ�Qׅr��2�e3���r+�4�j�
��?N1��(��!6߹�	ܝ�4%K8
���o4��2�`�=�m	�!&��a�!̔��G���A���Ll�$�:�4�Clb)\,4�X�7�F��d��t��1�:.%��~��~ktmP�T+k����(����5�J������ds�[��%t��+N{�I>�j6����J�A@�C�@=�jʒ^a��
��o��3�X�c��%�ʗ�Y�g��܇�i��UH�óu.UY[���M��R@�~c|�U�^X�]��<�D}X�t�5u��4�ǋ̢���W������jݐ��A�l��M�o'�av��^���mnuz;��}8��=��y�p`�)�o�k�,,�X�J]��/���k�c;?�l�FRN�h�1ꎈ%.fz��˅��nn�= �G��N�E������,Q�Rf}���+����7(n'�e��9���w���r����iwpU����d�Q��&}'i��`ǛÆ�~��g��A��4Ar��q?55du^�x^Y�xK�^�\]Z4��;׀ �hjV>��Є\+�W��0�0�FSzԒ�nQ,��g�5�5�� ^��7w@g�w������w�Cd��!���)��
�SOF��w�4��V�����)��VeA�J�d4T��e\*�T��UY49�w���M�������c��DuS{��ޱh8�$�Y�}^`��jј�H�a�y8�]����e����3	0�\E��$�p|򽠏����0 ^��9PJ��/xr}i�J��r=�i��O��a	�x,dm!sI�1Zܩ�����l�q��$�B�[���]����g;��̓��#;^�5Hr��0��tC\�l	'�s�t15�堔�z ���Xܰ��Վt�P�������S}���&f�!M�4!�r��'�P�����E�߼'Ω�'��݆�Q�^��E�R��)����w��JfI��b���Z��9PMJs( �سe���*�5�&C���/ɶ&����Q� W�I�G�&ka����`�gRc�jda�u�6 q6�jy̪
��fw�Z&t��ե =�A9#f1�s�y���l�C25��Ɓ���V�-��ͭ�@n�p,vhk�(ة���M���#���=.r,��zu�"�ࣧ���M&+��矞�tz5