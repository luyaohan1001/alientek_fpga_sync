// nios2os.v

// Generated using ACDS version 13.1 162 at 2019.01.29.15:19:08

`timescale 1 ps / 1 ps
module nios2os (
		input  wire        clk_clk,                    //            clk.clk
		input  wire        reset_reset_n,              //          reset.reset_n
		output wire [12:0] sdram_addr,                 //          sdram.addr
		output wire [1:0]  sdram_ba,                   //               .ba
		output wire        sdram_cas_n,                //               .cas_n
		output wire        sdram_cke,                  //               .cke
		output wire        sdram_cs_n,                 //               .cs_n
		inout  wire [15:0] sdram_dq,                   //               .dq
		output wire [1:0]  sdram_dqm,                  //               .dqm
		output wire        sdram_ras_n,                //               .ras_n
		output wire        sdram_we_n,                 //               .we_n
		output wire        epcs_flash_dclk,            //     epcs_flash.dclk
		output wire        epcs_flash_sce,             //               .sce
		output wire        epcs_flash_sdo,             //               .sdo
		input  wire        epcs_flash_data0,           //               .data0
		input  wire        tse_pcs_tx_clk_clk,         // tse_pcs_tx_clk.clk
		input  wire        tse_pcs_rx_clk_clk,         // tse_pcs_rx_clk.clk
		input  wire        tse_mac_stu_set_10,         //    tse_mac_stu.set_10
		input  wire        tse_mac_stu_set_1000,       //               .set_1000
		output wire        tse_mac_stu_eth_mode,       //               .eth_mode
		output wire        tse_mac_stu_ena_10,         //               .ena_10
		input  wire [3:0]  tse_mac_mii_rx_d,           //        tse_mac.mii_rx_d
		input  wire        tse_mac_mii_rx_dv,          //               .mii_rx_dv
		input  wire        tse_mac_mii_rx_err,         //               .mii_rx_err
		output wire [3:0]  tse_mac_mii_tx_d,           //               .mii_tx_d
		output wire        tse_mac_mii_tx_en,          //               .mii_tx_en
		output wire        tse_mac_mii_tx_err,         //               .mii_tx_err
		input  wire        tse_mac_misc_ff_tx_crc_fwd, //   tse_mac_misc.ff_tx_crc_fwd
		output wire        tse_mac_misc_ff_tx_septy,   //               .ff_tx_septy
		output wire        tse_mac_misc_tx_ff_uflow,   //               .tx_ff_uflow
		output wire        tse_mac_misc_ff_tx_a_full,  //               .ff_tx_a_full
		output wire        tse_mac_misc_ff_tx_a_empty, //               .ff_tx_a_empty
		output wire [17:0] tse_mac_misc_rx_err_stat,   //               .rx_err_stat
		output wire [3:0]  tse_mac_misc_rx_frm_type,   //               .rx_frm_type
		output wire        tse_mac_misc_ff_rx_dsav,    //               .ff_rx_dsav
		output wire        tse_mac_misc_ff_rx_a_full,  //               .ff_rx_a_full
		output wire        tse_mac_misc_ff_rx_a_empty, //               .ff_rx_a_empty
		output wire [3:0]  led_export                  //            led.export
	);

	wire         sgdma_tx_out_endofpacket;                                             // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire         sgdma_tx_out_valid;                                                   // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire         sgdma_tx_out_startofpacket;                                           // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire         sgdma_tx_out_error;                                                   // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                                   // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire  [31:0] sgdma_tx_out_data;                                                    // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire         sgdma_tx_out_ready;                                                   // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_writedata;                             // mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	wire   [3:0] mm_interconnect_0_sgdma_tx_csr_address;                               // mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	wire         mm_interconnect_0_sgdma_tx_csr_chipselect;                            // mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	wire         mm_interconnect_0_sgdma_tx_csr_write;                                 // mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	wire         mm_interconnect_0_sgdma_tx_csr_read;                                  // mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_readdata;                              // sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_writedata;                             // mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	wire   [3:0] mm_interconnect_0_sgdma_rx_csr_address;                               // mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	wire         mm_interconnect_0_sgdma_rx_csr_chipselect;                            // mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	wire         mm_interconnect_0_sgdma_rx_csr_write;                                 // mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	wire         mm_interconnect_0_sgdma_rx_csr_read;                                  // mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_readdata;                              // sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                   // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                  // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire         nios2_instruction_master_waitrequest;                                 // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [25:0] nios2_instruction_master_address;                                     // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                        // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                                    // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                               // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire  [31:0] mm_interconnect_0_descriptor_memory_s2_writedata;                     // mm_interconnect_0:descriptor_memory_s2_writedata -> descriptor_memory:writedata2
	wire   [6:0] mm_interconnect_0_descriptor_memory_s2_address;                       // mm_interconnect_0:descriptor_memory_s2_address -> descriptor_memory:address2
	wire         mm_interconnect_0_descriptor_memory_s2_chipselect;                    // mm_interconnect_0:descriptor_memory_s2_chipselect -> descriptor_memory:chipselect2
	wire         mm_interconnect_0_descriptor_memory_s2_clken;                         // mm_interconnect_0:descriptor_memory_s2_clken -> descriptor_memory:clken2
	wire         mm_interconnect_0_descriptor_memory_s2_write;                         // mm_interconnect_0:descriptor_memory_s2_write -> descriptor_memory:write2
	wire  [31:0] mm_interconnect_0_descriptor_memory_s2_readdata;                      // descriptor_memory:readdata2 -> mm_interconnect_0:descriptor_memory_s2_readdata
	wire   [3:0] mm_interconnect_0_descriptor_memory_s2_byteenable;                    // mm_interconnect_0:descriptor_memory_s2_byteenable -> descriptor_memory:byteenable2
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_controller_epcs_control_port_writedata -> epcs_flash_controller:writedata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_controller_epcs_control_port_address -> epcs_flash_controller:address
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_controller_epcs_control_port_chipselect -> epcs_flash_controller:chipselect
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_controller_epcs_control_port_write -> epcs_flash_controller:write_n
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_controller_epcs_control_port_read -> epcs_flash_controller:read_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata;   // epcs_flash_controller:readdata -> mm_interconnect_0:epcs_flash_controller_epcs_control_port_readdata
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_writedata;                        // mm_interconnect_0:high_res_timer_s1_writedata -> high_res_timer:writedata
	wire   [2:0] mm_interconnect_0_high_res_timer_s1_address;                          // mm_interconnect_0:high_res_timer_s1_address -> high_res_timer:address
	wire         mm_interconnect_0_high_res_timer_s1_chipselect;                       // mm_interconnect_0:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	wire         mm_interconnect_0_high_res_timer_s1_write;                            // mm_interconnect_0:high_res_timer_s1_write -> high_res_timer:write_n
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_readdata;                         // high_res_timer:readdata -> mm_interconnect_0:high_res_timer_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                               // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                 // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                   // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                     // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                      // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                  // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                             // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_tse_mac_control_port_waitrequest;                   // tse_mac:waitrequest -> mm_interconnect_0:tse_mac_control_port_waitrequest
	wire  [31:0] mm_interconnect_0_tse_mac_control_port_writedata;                     // mm_interconnect_0:tse_mac_control_port_writedata -> tse_mac:writedata
	wire   [7:0] mm_interconnect_0_tse_mac_control_port_address;                       // mm_interconnect_0:tse_mac_control_port_address -> tse_mac:address
	wire         mm_interconnect_0_tse_mac_control_port_write;                         // mm_interconnect_0:tse_mac_control_port_write -> tse_mac:write
	wire         mm_interconnect_0_tse_mac_control_port_read;                          // mm_interconnect_0:tse_mac_control_port_read -> tse_mac:read
	wire  [31:0] mm_interconnect_0_tse_mac_control_port_readdata;                      // tse_mac:readdata -> mm_interconnect_0:tse_mac_control_port_readdata
	wire         nios2_data_master_waitrequest;                                        // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                          // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [25:0] nios2_data_master_address;                                            // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                              // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                               // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                           // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                                        // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire         nios2_data_master_readdatavalid;                                      // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                                         // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;            // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;               // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                         // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                           // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                        // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                             // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                          // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;                // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;                  // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;                    // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;                      // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;                       // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;                   // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;                // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;                 // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;                               // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;                                 // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_0_led_pio_s1_chipselect;                              // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire         mm_interconnect_0_led_pio_s1_write;                                   // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;                                // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire   [0:0] pb_dma_to_sdram_m0_burstcount;                                        // pb_dma_to_sdram:m0_burstcount -> mm_interconnect_0:pb_dma_to_sdram_m0_burstcount
	wire         pb_dma_to_sdram_m0_waitrequest;                                       // mm_interconnect_0:pb_dma_to_sdram_m0_waitrequest -> pb_dma_to_sdram:m0_waitrequest
	wire  [26:0] pb_dma_to_sdram_m0_address;                                           // pb_dma_to_sdram:m0_address -> mm_interconnect_0:pb_dma_to_sdram_m0_address
	wire  [31:0] pb_dma_to_sdram_m0_writedata;                                         // pb_dma_to_sdram:m0_writedata -> mm_interconnect_0:pb_dma_to_sdram_m0_writedata
	wire         pb_dma_to_sdram_m0_write;                                             // pb_dma_to_sdram:m0_write -> mm_interconnect_0:pb_dma_to_sdram_m0_write
	wire         pb_dma_to_sdram_m0_read;                                              // pb_dma_to_sdram:m0_read -> mm_interconnect_0:pb_dma_to_sdram_m0_read
	wire  [31:0] pb_dma_to_sdram_m0_readdata;                                          // mm_interconnect_0:pb_dma_to_sdram_m0_readdata -> pb_dma_to_sdram:m0_readdata
	wire         pb_dma_to_sdram_m0_debugaccess;                                       // pb_dma_to_sdram:m0_debugaccess -> mm_interconnect_0:pb_dma_to_sdram_m0_debugaccess
	wire   [3:0] pb_dma_to_sdram_m0_byteenable;                                        // pb_dma_to_sdram:m0_byteenable -> mm_interconnect_0:pb_dma_to_sdram_m0_byteenable
	wire         pb_dma_to_sdram_m0_readdatavalid;                                     // mm_interconnect_0:pb_dma_to_sdram_m0_readdatavalid -> pb_dma_to_sdram:m0_readdatavalid
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_writedata;                     // mm_interconnect_1:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire   [6:0] mm_interconnect_1_descriptor_memory_s1_address;                       // mm_interconnect_1:descriptor_memory_s1_address -> descriptor_memory:address
	wire         mm_interconnect_1_descriptor_memory_s1_chipselect;                    // mm_interconnect_1:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire         mm_interconnect_1_descriptor_memory_s1_clken;                         // mm_interconnect_1:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_1_descriptor_memory_s1_write;                         // mm_interconnect_1:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_1_descriptor_memory_s1_readdata;                      // descriptor_memory:readdata -> mm_interconnect_1:descriptor_memory_s1_readdata
	wire   [3:0] mm_interconnect_1_descriptor_memory_s1_byteenable;                    // mm_interconnect_1:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         sgdma_tx_descriptor_write_waitrequest;                                // mm_interconnect_1:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                                  // sgdma_tx:descriptor_write_writedata -> mm_interconnect_1:sgdma_tx_descriptor_write_writedata
	wire  [31:0] sgdma_tx_descriptor_write_address;                                    // sgdma_tx:descriptor_write_address -> mm_interconnect_1:sgdma_tx_descriptor_write_address
	wire         sgdma_tx_descriptor_write_write;                                      // sgdma_tx:descriptor_write_write -> mm_interconnect_1:sgdma_tx_descriptor_write_write
	wire         sgdma_rx_descriptor_read_waitrequest;                                 // mm_interconnect_1:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                                     // sgdma_rx:descriptor_read_address -> mm_interconnect_1:sgdma_rx_descriptor_read_address
	wire         sgdma_rx_descriptor_read_read;                                        // sgdma_rx:descriptor_read_read -> mm_interconnect_1:sgdma_rx_descriptor_read_read
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                                    // mm_interconnect_1:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_readdatavalid;                               // mm_interconnect_1:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire         sgdma_tx_descriptor_read_waitrequest;                                 // mm_interconnect_1:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                                     // sgdma_tx:descriptor_read_address -> mm_interconnect_1:sgdma_tx_descriptor_read_address
	wire         sgdma_tx_descriptor_read_read;                                        // sgdma_tx:descriptor_read_read -> mm_interconnect_1:sgdma_tx_descriptor_read_read
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                                    // mm_interconnect_1:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_readdatavalid;                               // mm_interconnect_1:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire         sgdma_rx_descriptor_write_waitrequest;                                // mm_interconnect_1:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                                  // sgdma_rx:descriptor_write_writedata -> mm_interconnect_1:sgdma_rx_descriptor_write_writedata
	wire  [31:0] sgdma_rx_descriptor_write_address;                                    // sgdma_rx:descriptor_write_address -> mm_interconnect_1:sgdma_rx_descriptor_write_address
	wire         sgdma_rx_descriptor_write_write;                                      // sgdma_rx:descriptor_write_write -> mm_interconnect_1:sgdma_rx_descriptor_write_write
	wire         sgdma_tx_m_read_waitrequest;                                          // mm_interconnect_2:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                              // sgdma_tx:m_read_address -> mm_interconnect_2:sgdma_tx_m_read_address
	wire         sgdma_tx_m_read_read;                                                 // sgdma_tx:m_read_read -> mm_interconnect_2:sgdma_tx_m_read_read
	wire  [31:0] sgdma_tx_m_read_readdata;                                             // mm_interconnect_2:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_readdatavalid;                                        // mm_interconnect_2:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire         sgdma_rx_m_write_waitrequest;                                         // mm_interconnect_2:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_writedata;                                           // sgdma_rx:m_write_writedata -> mm_interconnect_2:sgdma_rx_m_write_writedata
	wire  [31:0] sgdma_rx_m_write_address;                                             // sgdma_rx:m_write_address -> mm_interconnect_2:sgdma_rx_m_write_address
	wire         sgdma_rx_m_write_write;                                               // sgdma_rx:m_write_write -> mm_interconnect_2:sgdma_rx_m_write_write
	wire   [3:0] sgdma_rx_m_write_byteenable;                                          // sgdma_rx:m_write_byteenable -> mm_interconnect_2:sgdma_rx_m_write_byteenable
	wire         mm_interconnect_2_pb_dma_to_sdram_s0_waitrequest;                     // pb_dma_to_sdram:s0_waitrequest -> mm_interconnect_2:pb_dma_to_sdram_s0_waitrequest
	wire   [0:0] mm_interconnect_2_pb_dma_to_sdram_s0_burstcount;                      // mm_interconnect_2:pb_dma_to_sdram_s0_burstcount -> pb_dma_to_sdram:s0_burstcount
	wire  [31:0] mm_interconnect_2_pb_dma_to_sdram_s0_writedata;                       // mm_interconnect_2:pb_dma_to_sdram_s0_writedata -> pb_dma_to_sdram:s0_writedata
	wire  [26:0] mm_interconnect_2_pb_dma_to_sdram_s0_address;                         // mm_interconnect_2:pb_dma_to_sdram_s0_address -> pb_dma_to_sdram:s0_address
	wire         mm_interconnect_2_pb_dma_to_sdram_s0_write;                           // mm_interconnect_2:pb_dma_to_sdram_s0_write -> pb_dma_to_sdram:s0_write
	wire         mm_interconnect_2_pb_dma_to_sdram_s0_read;                            // mm_interconnect_2:pb_dma_to_sdram_s0_read -> pb_dma_to_sdram:s0_read
	wire  [31:0] mm_interconnect_2_pb_dma_to_sdram_s0_readdata;                        // pb_dma_to_sdram:s0_readdata -> mm_interconnect_2:pb_dma_to_sdram_s0_readdata
	wire         mm_interconnect_2_pb_dma_to_sdram_s0_debugaccess;                     // mm_interconnect_2:pb_dma_to_sdram_s0_debugaccess -> pb_dma_to_sdram:s0_debugaccess
	wire         mm_interconnect_2_pb_dma_to_sdram_s0_readdatavalid;                   // pb_dma_to_sdram:s0_readdatavalid -> mm_interconnect_2:pb_dma_to_sdram_s0_readdatavalid
	wire   [3:0] mm_interconnect_2_pb_dma_to_sdram_s0_byteenable;                      // mm_interconnect_2:pb_dma_to_sdram_s0_byteenable -> pb_dma_to_sdram:s0_byteenable
	wire         irq_mapper_receiver0_irq;                                             // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                             // epcs_flash_controller:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                             // sgdma_tx:csr_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                             // sgdma_rx:csr_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                             // sys_clk_timer:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                             // high_res_timer:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_d_irq_irq;                                                      // irq_mapper:sender_irq -> nios2:d_irq
	wire         tse_mac_receive_endofpacket;                                          // tse_mac:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire         tse_mac_receive_valid;                                                // tse_mac:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire         tse_mac_receive_startofpacket;                                        // tse_mac:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire   [5:0] tse_mac_receive_error;                                                // tse_mac:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] tse_mac_receive_empty;                                                // tse_mac:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire  [31:0] tse_mac_receive_data;                                                 // tse_mac:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_mac_receive_ready;                                                // avalon_st_adapter:in_0_ready -> tse_mac:ff_rx_rdy
	wire         avalon_st_adapter_out_0_endofpacket;                                  // avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                        // avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	wire         avalon_st_adapter_out_0_startofpacket;                                // avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                                        // avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                                        // avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	wire  [31:0] avalon_st_adapter_out_0_data;                                         // avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	wire         avalon_st_adapter_out_0_ready;                                        // sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, descriptor_memory:reset2, epcs_flash_controller:reset_n, high_res_timer:reset_n, irq_mapper:reset, jtag_uart:rst_n, led_pio:reset_n, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:sgdma_rx_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sgdma_rx_reset_reset_bridge_in_reset_reset, nios2:reset_n, pb_dma_to_sdram:reset, rst_translator:in_reset, sdram:reset_n, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, sys_clk_timer:reset_n, sysid_qsys:reset_n, tse_mac:reset]
	wire         rst_controller_reset_out_reset_req;                                   // rst_controller:reset_req -> [descriptor_memory:reset_req, descriptor_memory:reset_req2, epcs_flash_controller:reset_req, nios2:reset_req, rst_translator:reset_req_in]
	wire         nios2_jtag_debug_module_reset_reset;                                  // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios2os_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	nios2os_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	nios2os_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	nios2os_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios2os_epcs_flash_controller epcs_flash_controller (
		.clk           (clk_clk),                                                              //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                      //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                                   //                  .reset_req
		.address       (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                                     //                  .dataavailable
		.endofpacket   (),                                                                     //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                                     //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver1_irq),                                             //               irq.irq
		.dclk          (epcs_flash_dclk),                                                      //          external.export
		.sce           (epcs_flash_sce),                                                       //                  .export
		.sdo           (epcs_flash_sdo),                                                       //                  .export
		.data0         (epcs_flash_data0)                                                      //                  .export
	);

	nios2os_tse_mac tse_mac (
		.clk           (clk_clk),                                            // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                     //              reset_connection.reset
		.address       (mm_interconnect_0_tse_mac_control_port_address),     //                  control_port.address
		.readdata      (mm_interconnect_0_tse_mac_control_port_readdata),    //                              .readdata
		.read          (mm_interconnect_0_tse_mac_control_port_read),        //                              .read
		.writedata     (mm_interconnect_0_tse_mac_control_port_writedata),   //                              .writedata
		.write         (mm_interconnect_0_tse_mac_control_port_write),       //                              .write
		.waitrequest   (mm_interconnect_0_tse_mac_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (tse_pcs_tx_clk_clk),                                 //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (tse_pcs_rx_clk_clk),                                 //   pcs_mac_rx_clock_connection.clk
		.set_10        (tse_mac_stu_set_10),                                 //         mac_status_connection.set_10
		.set_1000      (tse_mac_stu_set_1000),                               //                              .set_1000
		.eth_mode      (tse_mac_stu_eth_mode),                               //                              .eth_mode
		.ena_10        (tse_mac_stu_ena_10),                                 //                              .ena_10
		.m_rx_d        (tse_mac_mii_rx_d),                                   //            mac_mii_connection.mii_rx_d
		.m_rx_en       (tse_mac_mii_rx_dv),                                  //                              .mii_rx_dv
		.m_rx_err      (tse_mac_mii_rx_err),                                 //                              .mii_rx_err
		.m_tx_d        (tse_mac_mii_tx_d),                                   //                              .mii_tx_d
		.m_tx_en       (tse_mac_mii_tx_en),                                  //                              .mii_tx_en
		.m_tx_err      (tse_mac_mii_tx_err),                                 //                              .mii_tx_err
		.ff_rx_clk     (clk_clk),                                            //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                            //     transmit_clock_connection.clk
		.ff_rx_data    (tse_mac_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_mac_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_mac_receive_error),                              //                              .error
		.ff_rx_mod     (tse_mac_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_mac_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_mac_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_mac_receive_valid),                              //                              .valid
		.ff_tx_data    (sgdma_tx_out_data),                                  //                      transmit.data
		.ff_tx_eop     (sgdma_tx_out_endofpacket),                           //                              .endofpacket
		.ff_tx_err     (sgdma_tx_out_error),                                 //                              .error
		.ff_tx_mod     (sgdma_tx_out_empty),                                 //                              .empty
		.ff_tx_rdy     (sgdma_tx_out_ready),                                 //                              .ready
		.ff_tx_sop     (sgdma_tx_out_startofpacket),                         //                              .startofpacket
		.ff_tx_wren    (sgdma_tx_out_valid),                                 //                              .valid
		.ff_tx_crc_fwd (tse_mac_misc_ff_tx_crc_fwd),                         //           mac_misc_connection.ff_tx_crc_fwd
		.ff_tx_septy   (tse_mac_misc_ff_tx_septy),                           //                              .ff_tx_septy
		.tx_ff_uflow   (tse_mac_misc_tx_ff_uflow),                           //                              .tx_ff_uflow
		.ff_tx_a_full  (tse_mac_misc_ff_tx_a_full),                          //                              .ff_tx_a_full
		.ff_tx_a_empty (tse_mac_misc_ff_tx_a_empty),                         //                              .ff_tx_a_empty
		.rx_err_stat   (tse_mac_misc_rx_err_stat),                           //                              .rx_err_stat
		.rx_frm_type   (tse_mac_misc_rx_frm_type),                           //                              .rx_frm_type
		.ff_rx_dsav    (tse_mac_misc_ff_rx_dsav),                            //                              .ff_rx_dsav
		.ff_rx_a_full  (tse_mac_misc_ff_rx_a_full),                          //                              .ff_rx_a_full
		.ff_rx_a_empty (tse_mac_misc_ff_rx_a_empty)                          //                              .ff_rx_a_empty
	);

	nios2os_sgdma_tx sgdma_tx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_tx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_tx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_tx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_tx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_tx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_tx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver2_irq),                  //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                      //                 .read
		.out_data                      (sgdma_tx_out_data),                         //              out.data
		.out_valid                     (sgdma_tx_out_valid),                        //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                        //                 .empty
		.out_error                     (sgdma_tx_out_error)                         //                 .error
	);

	nios2os_sgdma_rx sgdma_rx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_rx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_rx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_rx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_rx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_rx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_rx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver3_irq),                  //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),     //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),       //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),              //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),             //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),             //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),             //                 .empty
		.in_error                      (avalon_st_adapter_out_0_error),             //                 .error
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable)                //                 .byteenable
	);

	nios2os_descriptor_memory descriptor_memory (
		.clk         (clk_clk),                                           //   clk1.clk
		.address     (mm_interconnect_1_descriptor_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_descriptor_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_descriptor_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_descriptor_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_1_descriptor_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_descriptor_memory_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                    // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),                //       .reset_req
		.address2    (mm_interconnect_0_descriptor_memory_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_descriptor_memory_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_descriptor_memory_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_descriptor_memory_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_descriptor_memory_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_descriptor_memory_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_descriptor_memory_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                           //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                    // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)                 //       .reset_req
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pb_dma_to_sdram (
		.clk              (clk_clk),                                            //   clk.clk
		.reset            (rst_controller_reset_out_reset),                     // reset.reset
		.s0_waitrequest   (mm_interconnect_2_pb_dma_to_sdram_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_2_pb_dma_to_sdram_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_2_pb_dma_to_sdram_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_2_pb_dma_to_sdram_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_2_pb_dma_to_sdram_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_2_pb_dma_to_sdram_s0_address),       //      .address
		.s0_write         (mm_interconnect_2_pb_dma_to_sdram_s0_write),         //      .write
		.s0_read          (mm_interconnect_2_pb_dma_to_sdram_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_2_pb_dma_to_sdram_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_2_pb_dma_to_sdram_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pb_dma_to_sdram_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pb_dma_to_sdram_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pb_dma_to_sdram_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pb_dma_to_sdram_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pb_dma_to_sdram_m0_writedata),                       //      .writedata
		.m0_address       (pb_dma_to_sdram_m0_address),                         //      .address
		.m0_write         (pb_dma_to_sdram_m0_write),                           //      .write
		.m0_read          (pb_dma_to_sdram_m0_read),                            //      .read
		.m0_byteenable    (pb_dma_to_sdram_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pb_dma_to_sdram_m0_debugaccess)                      //      .debugaccess
	);

	nios2os_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                       //   irq.irq
	);

	nios2os_high_res_timer high_res_timer (
		.clk        (clk_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_high_res_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                        //   irq.irq
	);

	nios2os_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_export)                               // external_connection.export
	);

	nios2os_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                        (clk_clk),                                                              //                                 clk_clk.clk
		.nios2_reset_n_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                                       //     nios2_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                          (nios2_data_master_address),                                            //                       nios2_data_master.address
		.nios2_data_master_waitrequest                      (nios2_data_master_waitrequest),                                        //                                        .waitrequest
		.nios2_data_master_byteenable                       (nios2_data_master_byteenable),                                         //                                        .byteenable
		.nios2_data_master_read                             (nios2_data_master_read),                                               //                                        .read
		.nios2_data_master_readdata                         (nios2_data_master_readdata),                                           //                                        .readdata
		.nios2_data_master_readdatavalid                    (nios2_data_master_readdatavalid),                                      //                                        .readdatavalid
		.nios2_data_master_write                            (nios2_data_master_write),                                              //                                        .write
		.nios2_data_master_writedata                        (nios2_data_master_writedata),                                          //                                        .writedata
		.nios2_data_master_debugaccess                      (nios2_data_master_debugaccess),                                        //                                        .debugaccess
		.nios2_instruction_master_address                   (nios2_instruction_master_address),                                     //                nios2_instruction_master.address
		.nios2_instruction_master_waitrequest               (nios2_instruction_master_waitrequest),                                 //                                        .waitrequest
		.nios2_instruction_master_read                      (nios2_instruction_master_read),                                        //                                        .read
		.nios2_instruction_master_readdata                  (nios2_instruction_master_readdata),                                    //                                        .readdata
		.nios2_instruction_master_readdatavalid             (nios2_instruction_master_readdatavalid),                               //                                        .readdatavalid
		.pb_dma_to_sdram_m0_address                         (pb_dma_to_sdram_m0_address),                                           //                      pb_dma_to_sdram_m0.address
		.pb_dma_to_sdram_m0_waitrequest                     (pb_dma_to_sdram_m0_waitrequest),                                       //                                        .waitrequest
		.pb_dma_to_sdram_m0_burstcount                      (pb_dma_to_sdram_m0_burstcount),                                        //                                        .burstcount
		.pb_dma_to_sdram_m0_byteenable                      (pb_dma_to_sdram_m0_byteenable),                                        //                                        .byteenable
		.pb_dma_to_sdram_m0_read                            (pb_dma_to_sdram_m0_read),                                              //                                        .read
		.pb_dma_to_sdram_m0_readdata                        (pb_dma_to_sdram_m0_readdata),                                          //                                        .readdata
		.pb_dma_to_sdram_m0_readdatavalid                   (pb_dma_to_sdram_m0_readdatavalid),                                     //                                        .readdatavalid
		.pb_dma_to_sdram_m0_write                           (pb_dma_to_sdram_m0_write),                                             //                                        .write
		.pb_dma_to_sdram_m0_writedata                       (pb_dma_to_sdram_m0_writedata),                                         //                                        .writedata
		.pb_dma_to_sdram_m0_debugaccess                     (pb_dma_to_sdram_m0_debugaccess),                                       //                                        .debugaccess
		.descriptor_memory_s2_address                       (mm_interconnect_0_descriptor_memory_s2_address),                       //                    descriptor_memory_s2.address
		.descriptor_memory_s2_write                         (mm_interconnect_0_descriptor_memory_s2_write),                         //                                        .write
		.descriptor_memory_s2_readdata                      (mm_interconnect_0_descriptor_memory_s2_readdata),                      //                                        .readdata
		.descriptor_memory_s2_writedata                     (mm_interconnect_0_descriptor_memory_s2_writedata),                     //                                        .writedata
		.descriptor_memory_s2_byteenable                    (mm_interconnect_0_descriptor_memory_s2_byteenable),                    //                                        .byteenable
		.descriptor_memory_s2_chipselect                    (mm_interconnect_0_descriptor_memory_s2_chipselect),                    //                                        .chipselect
		.descriptor_memory_s2_clken                         (mm_interconnect_0_descriptor_memory_s2_clken),                         //                                        .clken
		.epcs_flash_controller_epcs_control_port_address    (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    // epcs_flash_controller_epcs_control_port.address
		.epcs_flash_controller_epcs_control_port_write      (mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),      //                                        .write
		.epcs_flash_controller_epcs_control_port_read       (mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),       //                                        .read
		.epcs_flash_controller_epcs_control_port_readdata   (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                                        .readdata
		.epcs_flash_controller_epcs_control_port_writedata  (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                                        .writedata
		.epcs_flash_controller_epcs_control_port_chipselect (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                                        .chipselect
		.high_res_timer_s1_address                          (mm_interconnect_0_high_res_timer_s1_address),                          //                       high_res_timer_s1.address
		.high_res_timer_s1_write                            (mm_interconnect_0_high_res_timer_s1_write),                            //                                        .write
		.high_res_timer_s1_readdata                         (mm_interconnect_0_high_res_timer_s1_readdata),                         //                                        .readdata
		.high_res_timer_s1_writedata                        (mm_interconnect_0_high_res_timer_s1_writedata),                        //                                        .writedata
		.high_res_timer_s1_chipselect                       (mm_interconnect_0_high_res_timer_s1_chipselect),                       //                                        .chipselect
		.jtag_uart_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                //             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                  //                                        .write
		.jtag_uart_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                   //                                        .read
		.jtag_uart_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),               //                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),              //                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),            //                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),             //                                        .chipselect
		.led_pio_s1_address                                 (mm_interconnect_0_led_pio_s1_address),                                 //                              led_pio_s1.address
		.led_pio_s1_write                                   (mm_interconnect_0_led_pio_s1_write),                                   //                                        .write
		.led_pio_s1_readdata                                (mm_interconnect_0_led_pio_s1_readdata),                                //                                        .readdata
		.led_pio_s1_writedata                               (mm_interconnect_0_led_pio_s1_writedata),                               //                                        .writedata
		.led_pio_s1_chipselect                              (mm_interconnect_0_led_pio_s1_chipselect),                              //                                        .chipselect
		.nios2_jtag_debug_module_address                    (mm_interconnect_0_nios2_jtag_debug_module_address),                    //                 nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write                      (mm_interconnect_0_nios2_jtag_debug_module_write),                      //                                        .write
		.nios2_jtag_debug_module_read                       (mm_interconnect_0_nios2_jtag_debug_module_read),                       //                                        .read
		.nios2_jtag_debug_module_readdata                   (mm_interconnect_0_nios2_jtag_debug_module_readdata),                   //                                        .readdata
		.nios2_jtag_debug_module_writedata                  (mm_interconnect_0_nios2_jtag_debug_module_writedata),                  //                                        .writedata
		.nios2_jtag_debug_module_byteenable                 (mm_interconnect_0_nios2_jtag_debug_module_byteenable),                 //                                        .byteenable
		.nios2_jtag_debug_module_waitrequest                (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),                //                                        .waitrequest
		.nios2_jtag_debug_module_debugaccess                (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),                //                                        .debugaccess
		.sdram_s1_address                                   (mm_interconnect_0_sdram_s1_address),                                   //                                sdram_s1.address
		.sdram_s1_write                                     (mm_interconnect_0_sdram_s1_write),                                     //                                        .write
		.sdram_s1_read                                      (mm_interconnect_0_sdram_s1_read),                                      //                                        .read
		.sdram_s1_readdata                                  (mm_interconnect_0_sdram_s1_readdata),                                  //                                        .readdata
		.sdram_s1_writedata                                 (mm_interconnect_0_sdram_s1_writedata),                                 //                                        .writedata
		.sdram_s1_byteenable                                (mm_interconnect_0_sdram_s1_byteenable),                                //                                        .byteenable
		.sdram_s1_readdatavalid                             (mm_interconnect_0_sdram_s1_readdatavalid),                             //                                        .readdatavalid
		.sdram_s1_waitrequest                               (mm_interconnect_0_sdram_s1_waitrequest),                               //                                        .waitrequest
		.sdram_s1_chipselect                                (mm_interconnect_0_sdram_s1_chipselect),                                //                                        .chipselect
		.sgdma_rx_csr_address                               (mm_interconnect_0_sgdma_rx_csr_address),                               //                            sgdma_rx_csr.address
		.sgdma_rx_csr_write                                 (mm_interconnect_0_sgdma_rx_csr_write),                                 //                                        .write
		.sgdma_rx_csr_read                                  (mm_interconnect_0_sgdma_rx_csr_read),                                  //                                        .read
		.sgdma_rx_csr_readdata                              (mm_interconnect_0_sgdma_rx_csr_readdata),                              //                                        .readdata
		.sgdma_rx_csr_writedata                             (mm_interconnect_0_sgdma_rx_csr_writedata),                             //                                        .writedata
		.sgdma_rx_csr_chipselect                            (mm_interconnect_0_sgdma_rx_csr_chipselect),                            //                                        .chipselect
		.sgdma_tx_csr_address                               (mm_interconnect_0_sgdma_tx_csr_address),                               //                            sgdma_tx_csr.address
		.sgdma_tx_csr_write                                 (mm_interconnect_0_sgdma_tx_csr_write),                                 //                                        .write
		.sgdma_tx_csr_read                                  (mm_interconnect_0_sgdma_tx_csr_read),                                  //                                        .read
		.sgdma_tx_csr_readdata                              (mm_interconnect_0_sgdma_tx_csr_readdata),                              //                                        .readdata
		.sgdma_tx_csr_writedata                             (mm_interconnect_0_sgdma_tx_csr_writedata),                             //                                        .writedata
		.sgdma_tx_csr_chipselect                            (mm_interconnect_0_sgdma_tx_csr_chipselect),                            //                                        .chipselect
		.sys_clk_timer_s1_address                           (mm_interconnect_0_sys_clk_timer_s1_address),                           //                        sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                             (mm_interconnect_0_sys_clk_timer_s1_write),                             //                                        .write
		.sys_clk_timer_s1_readdata                          (mm_interconnect_0_sys_clk_timer_s1_readdata),                          //                                        .readdata
		.sys_clk_timer_s1_writedata                         (mm_interconnect_0_sys_clk_timer_s1_writedata),                         //                                        .writedata
		.sys_clk_timer_s1_chipselect                        (mm_interconnect_0_sys_clk_timer_s1_chipselect),                        //                                        .chipselect
		.sysid_qsys_control_slave_address                   (mm_interconnect_0_sysid_qsys_control_slave_address),                   //                sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                  (mm_interconnect_0_sysid_qsys_control_slave_readdata),                  //                                        .readdata
		.tse_mac_control_port_address                       (mm_interconnect_0_tse_mac_control_port_address),                       //                    tse_mac_control_port.address
		.tse_mac_control_port_write                         (mm_interconnect_0_tse_mac_control_port_write),                         //                                        .write
		.tse_mac_control_port_read                          (mm_interconnect_0_tse_mac_control_port_read),                          //                                        .read
		.tse_mac_control_port_readdata                      (mm_interconnect_0_tse_mac_control_port_readdata),                      //                                        .readdata
		.tse_mac_control_port_writedata                     (mm_interconnect_0_tse_mac_control_port_writedata),                     //                                        .writedata
		.tse_mac_control_port_waitrequest                   (mm_interconnect_0_tse_mac_control_port_waitrequest)                    //                                        .waitrequest
	);

	nios2os_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                                (clk_clk),                                           //                              clk_clk.clk
		.sgdma_rx_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // sgdma_rx_reset_reset_bridge_in_reset.reset
		.sgdma_rx_descriptor_read_address           (sgdma_rx_descriptor_read_address),                  //             sgdma_rx_descriptor_read.address
		.sgdma_rx_descriptor_read_waitrequest       (sgdma_rx_descriptor_read_waitrequest),              //                                     .waitrequest
		.sgdma_rx_descriptor_read_read              (sgdma_rx_descriptor_read_read),                     //                                     .read
		.sgdma_rx_descriptor_read_readdata          (sgdma_rx_descriptor_read_readdata),                 //                                     .readdata
		.sgdma_rx_descriptor_read_readdatavalid     (sgdma_rx_descriptor_read_readdatavalid),            //                                     .readdatavalid
		.sgdma_rx_descriptor_write_address          (sgdma_rx_descriptor_write_address),                 //            sgdma_rx_descriptor_write.address
		.sgdma_rx_descriptor_write_waitrequest      (sgdma_rx_descriptor_write_waitrequest),             //                                     .waitrequest
		.sgdma_rx_descriptor_write_write            (sgdma_rx_descriptor_write_write),                   //                                     .write
		.sgdma_rx_descriptor_write_writedata        (sgdma_rx_descriptor_write_writedata),               //                                     .writedata
		.sgdma_tx_descriptor_read_address           (sgdma_tx_descriptor_read_address),                  //             sgdma_tx_descriptor_read.address
		.sgdma_tx_descriptor_read_waitrequest       (sgdma_tx_descriptor_read_waitrequest),              //                                     .waitrequest
		.sgdma_tx_descriptor_read_read              (sgdma_tx_descriptor_read_read),                     //                                     .read
		.sgdma_tx_descriptor_read_readdata          (sgdma_tx_descriptor_read_readdata),                 //                                     .readdata
		.sgdma_tx_descriptor_read_readdatavalid     (sgdma_tx_descriptor_read_readdatavalid),            //                                     .readdatavalid
		.sgdma_tx_descriptor_write_address          (sgdma_tx_descriptor_write_address),                 //            sgdma_tx_descriptor_write.address
		.sgdma_tx_descriptor_write_waitrequest      (sgdma_tx_descriptor_write_waitrequest),             //                                     .waitrequest
		.sgdma_tx_descriptor_write_write            (sgdma_tx_descriptor_write_write),                   //                                     .write
		.sgdma_tx_descriptor_write_writedata        (sgdma_tx_descriptor_write_writedata),               //                                     .writedata
		.descriptor_memory_s1_address               (mm_interconnect_1_descriptor_memory_s1_address),    //                 descriptor_memory_s1.address
		.descriptor_memory_s1_write                 (mm_interconnect_1_descriptor_memory_s1_write),      //                                     .write
		.descriptor_memory_s1_readdata              (mm_interconnect_1_descriptor_memory_s1_readdata),   //                                     .readdata
		.descriptor_memory_s1_writedata             (mm_interconnect_1_descriptor_memory_s1_writedata),  //                                     .writedata
		.descriptor_memory_s1_byteenable            (mm_interconnect_1_descriptor_memory_s1_byteenable), //                                     .byteenable
		.descriptor_memory_s1_chipselect            (mm_interconnect_1_descriptor_memory_s1_chipselect), //                                     .chipselect
		.descriptor_memory_s1_clken                 (mm_interconnect_1_descriptor_memory_s1_clken)       //                                     .clken
	);

	nios2os_mm_interconnect_2 mm_interconnect_2 (
		.clk_clk_clk                                (clk_clk),                                            //                              clk_clk.clk
		.sgdma_rx_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // sgdma_rx_reset_reset_bridge_in_reset.reset
		.sgdma_rx_m_write_address                   (sgdma_rx_m_write_address),                           //                     sgdma_rx_m_write.address
		.sgdma_rx_m_write_waitrequest               (sgdma_rx_m_write_waitrequest),                       //                                     .waitrequest
		.sgdma_rx_m_write_byteenable                (sgdma_rx_m_write_byteenable),                        //                                     .byteenable
		.sgdma_rx_m_write_write                     (sgdma_rx_m_write_write),                             //                                     .write
		.sgdma_rx_m_write_writedata                 (sgdma_rx_m_write_writedata),                         //                                     .writedata
		.sgdma_tx_m_read_address                    (sgdma_tx_m_read_address),                            //                      sgdma_tx_m_read.address
		.sgdma_tx_m_read_waitrequest                (sgdma_tx_m_read_waitrequest),                        //                                     .waitrequest
		.sgdma_tx_m_read_read                       (sgdma_tx_m_read_read),                               //                                     .read
		.sgdma_tx_m_read_readdata                   (sgdma_tx_m_read_readdata),                           //                                     .readdata
		.sgdma_tx_m_read_readdatavalid              (sgdma_tx_m_read_readdatavalid),                      //                                     .readdatavalid
		.pb_dma_to_sdram_s0_address                 (mm_interconnect_2_pb_dma_to_sdram_s0_address),       //                   pb_dma_to_sdram_s0.address
		.pb_dma_to_sdram_s0_write                   (mm_interconnect_2_pb_dma_to_sdram_s0_write),         //                                     .write
		.pb_dma_to_sdram_s0_read                    (mm_interconnect_2_pb_dma_to_sdram_s0_read),          //                                     .read
		.pb_dma_to_sdram_s0_readdata                (mm_interconnect_2_pb_dma_to_sdram_s0_readdata),      //                                     .readdata
		.pb_dma_to_sdram_s0_writedata               (mm_interconnect_2_pb_dma_to_sdram_s0_writedata),     //                                     .writedata
		.pb_dma_to_sdram_s0_burstcount              (mm_interconnect_2_pb_dma_to_sdram_s0_burstcount),    //                                     .burstcount
		.pb_dma_to_sdram_s0_byteenable              (mm_interconnect_2_pb_dma_to_sdram_s0_byteenable),    //                                     .byteenable
		.pb_dma_to_sdram_s0_readdatavalid           (mm_interconnect_2_pb_dma_to_sdram_s0_readdatavalid), //                                     .readdatavalid
		.pb_dma_to_sdram_s0_waitrequest             (mm_interconnect_2_pb_dma_to_sdram_s0_waitrequest),   //                                     .waitrequest
		.pb_dma_to_sdram_s0_debugaccess             (mm_interconnect_2_pb_dma_to_sdram_s0_debugaccess)    //                                     .debugaccess
	);

	nios2os_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	nios2os_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_ready          (tse_mac_receive_ready),                 //     in_0.ready
		.in_0_valid          (tse_mac_receive_valid),                 //         .valid
		.in_0_data           (tse_mac_receive_data),                  //         .data
		.in_0_startofpacket  (tse_mac_receive_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (tse_mac_receive_endofpacket),           //         .endofpacket
		.in_0_empty          (tse_mac_receive_empty),                 //         .empty
		.in_0_error          (tse_mac_receive_error),                 //         .error
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //    out_0.ready
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_data          (avalon_st_adapter_out_0_data),          //         .data
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
