��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��>��@K�gP�Iuz�8n�?"1_����1&O��]���>qKw�#�\t����P��X�¿�_]�e���B*�-~�K��F��	b��Ī�46�b=ӛ+An��g�, 9���a��ID�es��lc�"���?Ef�����{MQ%��T��waoK�l�	d-O�8^F�g����+ZEʗ�5Ɉ�_�bV�~������оdP��S�����%������;�FotT����wx�c�av?��q���0��t�e9�K)�$]n��Q�k�ڸ� gwڸv��PnG$bj�u��%�3~� �L88��D	�9rX��.�v��6�K�Ȇa_j�kW�洊bH�0�?H�hg�ZvZKR崆vC0lңr�v�;�f�{Fi�>蛑9J���T>i��2�`���J=W�J*?MR#=����i�����7���p�+v�]}����%��u���>�@P�`��({�(��a��/}g��,��WF�HY�(��p�:�%P>ZP-\d�U̾�Np�9R^�<�'|����!������w/7�5��%�k��[��k����D^S��U!s�ǙoCM��>	X��1~`���rM6��[iZH�B| ��v�٩O�8�o�9T]r�T���H�1�zS|�b���O��K�����
��#|򐗪�$n[�s�p����f'�,���ސ�ÙS��=Ý��z�� �i�zY�_��,���dD����y{x�w��Z���N�Hd�w�R9��|`��h��^����fy�	�l�R�D/���@bf�Ÿ�iR
�Q�QEw�GS���4���$�h�Ϝ�R�[����'���<���gi�_��,GS�����4^�nY�Y��N�������ɢШUw.\�M�(y±˪4E���}���?���_
j@��S!���9��ř���p����#����������>h��P�}KK��7�ao�.|�iX�*U8 �����T����V,�s��O���,����O0i�l�ΧjZ��+Ş�%���d(�<&�]�^�p�[��&�{�L'?��$��oa�e��+#�|I�Na�/6<��R�p�|GL��RY-�#H4n���ݺse���@�e��՗�A1(��y���y���rT5�d�1U������tM�cQ/������s/1f>@���v���;o�FD$%��E I6S��{t;�k�X�M#bn��Ob��T�7!B%{�/�&F-��'������K����� =����Ais��Z�Sq9�H�v�/��1y����xU�YV�޹�^T���6�U9:�s��
�lҢ���$_������{_O��:��̬5m�컠{����g����#�B5g�����̃o�}�yc��C��9&���iK���X�[$�����Qi��pI9j�A��&Cfٛ�<J����HЮ)c�e�k�
`�b(�fQ�O�/j��H�\�z��˱��CQ�&74Õ� f F��I�A�Uztcǻ";��^��YW�x���<��]���*�%|��S9�G��(��И7��폌g����� -�Sٗ�6�wر�ߓ`{騞}��%ns�[lf����|-�P%�<��Ҩp�,>tFK���]*=9���&�c���M��:�w���7d�Q� �1[\]B�t��d�o���ʘ��)��j?��BAܖ yCl'�ͣ�Zp�����5,H,g��H���o"�(5F��i���aP������nŕ��ʺ%-���X����V��1�:���~0弪�?|��n�x��R��L���鵒o%K��B����]R0d��ݍf
�e��-�~�����G�ݻ��1�6�<�Qn�9ú���R��c�,�v�A�kr��k�J>�S��l�U����@�D��%����=o�\��#`�Ό4K�s�@�Q��]�{z5z��\;�<E�#�.{��A���-J�����!���>ǧ�a�5�W{]��*�r#�c����V3c��S�+��.�ƕ����']cF�7N����!�D�A���.���?k�t^�\��7���.�?2�X��9�W���t�]�੥��A2���*k\��?j�I�ɍ�C�l�ǹ�({��:�h���2i��i��F�?kO�~a�3�4�X�l��d�|�,ɨ:�����_�R���xm��l�G�7b�^�P .�蕄��`�����?�Ac�@�Ir���a��2	��{X�Pk�4�VJ��IW	�Z���As�$w�E��܋�R��ǿ0\	ùX��gIK�l�r�:���jJ.�t�sB�Q��3d��%dՅCP�rGi��1����6�g�