��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�^͉�������L�"�4�RW�������&������l�d9l�Gv�`.�0����N�P������b)���cڬ��kuK��"�5�&���w
UA�2ޭIɡv,h���
�>�����X�d�*<������F��h.]�{�W\�=^����k׵[�(�Ui��[.1���Bx�]��ٯH�ө�2���K��������(	�Y?DyE��/�
�k�U�Sߢ�h]��*i�C�� 6$�΅T� 3�տcf���-VpZlT���Le��e·���������F�\�ЗW��z��m�횖���$�x ��j��-Za9�!��0�����̛S���� N��SbZ-GWc�T�y$�[���9��k�>*��w x � $�D�7��~��ο�B�[��=����� T����B~��"\-Jgy��͇=�[��2�^�x��-�y��(���S���.G��+��oL?T�9�$�4]WD�n�Q���s��c�ܚ�����Gꚇ)���J�wZ���3uw�D�|��ԯ�C� e�o��]��x��o>R/%��n��ۡ��{xQ�J6�.>,�m!'�s��<�5���oTm1IՌ���[q�n.�O� =��H��9� @��,p�]���Kw��ϐ6+�r���9�Sı����4G�$��������A�@C�>�
���BAN����?��H������R3�@�w@�R(����Y����nW�-����':��'u�A�r��rs.[�N0�z!˽c�g���&ݜE�{�V_��Gw�o�lb�O�����]�@)x ����/��QH/屴�P�@���e�J�g��{��?)�S�Z��K�	���jfOG��Yg%ߞk����DY71Z��'tYv/�,G�~M���ڐPP��V�@�=��
2
GT!���M/�T-���OW�({2�:���������tU޶6�X���y��(A����U̺6�.�N�����t$<��O��Wܿ�s`GR^��Y5����T����e6yf1��v ���O�����G��:FK��Aom˔,܊���	�6���D�i���Z^��7r��U��.��MHE�?�U�]�Y�\{�����/���	�Y�O�Ҹ���^v|��d.�)0��l�h;���˟��a+q}�����C|��m2�#� DL/���÷P�/H�+��_<q @2��T�Jb�n�~�"*$S�篂DA�Y@[���*�<�2tn�l��|���u!ˀMC ��N�W.�l�ٌS�-�Q��;y_7���&Q0f#\�B��&q�7�i�PF��~m����-����Qt�O�vG���̐�J���a��b�������|�V��$��!�DiT��l+r��$z��"�۱y ���G��K����A�m�P��N���`8�T
3�R��q7��	�����r�����Q�� (�a��GO|oDS��lc�1ś�X����Oļ��řhUw�$CC"=��t���G��H�DY��A�m��b�!	�3[
��N��/��R�Q��jm:���&[�����flY��/�ܞ���lP�L�4��Di�.	������v�G�+�\��Ѣ+N�{�4�_g�T�����X��8u�蛣�.�)�� w0�"|�$��~}(��s�e<G|�M�?s����1�r<�&�V����u��v_A�X_5����p;��@+o6-��� ��m�� ��U�-P2�0���j�
<}��L�d��!=�N�۹�2^/7 b����۹f@��S����Y�*��&|�a�-�f�J��Gf)��`�Ή9
�������|�l���ʉiu�}-��ʝ
I��P�{�D� �7W@������uc"�!H�Y�4|5@��jPQ���9�œ��7Eߗ�{��"3�h���*��^��y���o/�,ܩ�=�j7n!SpI*�������ٳ)E8ǌ2�����ҹ6���6�
�J�l-C�%Pz�P����Qi䪿7���L�ɾqcp�^�s@��	N�@�b��z��0Z��>�n�F+�{�4��8���B����d-bz�(�����_St	��A��gjx0�C�$֙����XP��x�z�f҉Hշ�b
�&�A��oolݭJ#0�n�D���e^:�e�gn������ PcL�UQj���X���%�Ҥh]�=a�ϰ�e�Z���1�@�Πi#Z�i�j�]to�����T4�q|EBO�rv�/V��q~v���h���PF����;�̓�!9G���|�t����
r!����e��V鑧N�V'��˯<1��Z;��-m]�ؘ;�E5��i�OɠvJ���8T���H|���S�r�4Y���!R2�L�\I����a{��KWB�Y�"�ӻe'�\7x���Y�'�mM�!�q~R�sY���n7�1Е����-�c���Os��j�G:yj%z����Q�Ҩr����TT[37ӣB�2�V]���ȼ���Ɵ���?BvJ�p=��oF����x)�K���wo�m������N4���f���Q����|��~��ȷd��ʃ�A�����k�+G�}�����a�)�ahd�ሎ,���4d�}߈Q,$�=wP���?�	�#]%���IL���r�U$��r�Qq�sJI��;W��И����j�W���$�{=���"�Ե����������%�R9�!�lq�����z�ZG!L�eT��鈫�U����k�x=q�/_]�kc�$�!D�!3�$qv�'ߦ��F��e�.������DDx���!��i7��gkL�
s@������\���R�w�҆wb��nm\�8�J	ܣ%j�磍����׾�5�i���D�N���Wp�q�[���]�]��E$(9^�)ٲ��1�#~�{��hN��w�[p��\��>n��W�%PeFW�c�df&4�푭�e֌ ����ۚ�Wlp6�q'��o��C:n$�jq���U747Zv���h-4dx&`]��1/�{�8�.�P>'��b�(
��j�ِ�ά�� &��3����1ּ� xJ�9��]g���=!@��%�Ɔw\�
�� C��U��F����w�#�w�͗旧#45��Ru#��(HpJ�U`Kϥ�Q/V�zEه�L~-$�f�a����.!��HCU�G tS�U�ɬ�,]������Pc㳏IKhfU˽6�f����i(�yC���2�o�c�8��*�\�ƅ1��:�a�����8O^<T��Ô��j��*��㏢�I�@��]�-���'���%q?\�g{tN0vunG� l�����bΆe���=������C.R�jA�d���l�'�y�7��ov����M�܊ep�r0��rF�G�ly�h5�*L���YbH�~AK�ӕ�x�!.׬�tqB
=��s��l����0�=3Q�q�y�%#��ڽ��8!^P��F�9W%q�bz�)��_4�@�J-!�IM/0:��ď��4�XP��Y�/��V��@�f
��b���̸UU��Y��r�my3|��0���/����c	��,��c��T!��iV2>�����T��J����~�v��/]��>��#�S�����#��+�j����'�Ʒ�I^��ݧof���_�%�,�K���gwUx�Pae�����6�J���F��ڴ~�b �xJ�%Y=Z�J�z�Q������iޑ�W���&�k��
�&_���:I�C^����y�1]*��y���#��5�����\/q����i�D���o�B��2�`,�������O�hb��L}6��q4
�m�Sy�ȑ*֫�aȩː�4��(�W���:�����_�� |��J��;��&�o��#�Ԣ�L�	S����aԕ�%c�&)\3�6fHW_'m����h�RS����0O�M����Ӑ���=d����jo��9Jǎ�|�������Z(`(N�$�b��x��������z(�:��Ӄ%1�X&�w�R)z��Ho�W׎�B9AC����6"�h��@����w��!�XK�6�j����lC&��a�2[O��K�������^Er�xD��TC@<o� ��2�����}��m���J�5�Ѷ�b�ǻ�K��6�#
��S�����
[��%��]�\껁 յ�I��q�j`�hk�4���ϡ}Rn����dD������}�֞@a�8�V���qg���͠ж�� �W�����>-1J�]�p^z�9j��V,/��Z���--�ivj��O�(�A�F�{!v�)8
�c�Q�#C��ԍY�@;t@� ���1����qx����FW�c���m��T��8H���N��SPjPc���P��u��1��X�����d�:H��D�:J�W?v?ğ��#iu������ͮ�l���ݮ1�����\ꩌP�|]�P�ALU�Pȱl�����.>�]8a۹��y�c���B.�i�ډ'�[�b��F��E��5�b�XZ�
=��O�[|�����nXqtg��m%#������=A�@�V}3��)������v/#����D7�RsJ|��� ���9n��k�?�[�j������K,Ĺ~������Svb̩cl�x�4���5r��2B���f��1��sS����8� *��z�Lɧ���fL�ьn��)�T#2B�}�H�q�~j���g�)���1��<��q۞C����\����f�Z��U���6S��쒯��X8��W%,�B��q�4d `�Wrw�� ��~pG7*X��c��l�Tx�)!�����Tj�/�2���2oo�0�c��P�����Л�\,Dֈn�P����Q����4!;;�3X�O9WG�����>�����R>�V�,��.��GE5�:� QP!�D܄���+ щR�&n�X�s��B��)���2�L��t�[�x���L�p�[���Pdn��]`��Sh.�wg���,on0pU�+-Dg�����m9x���=g=x�\�C2c�BV�C�tY6v��g0LE�J# � �c�zTv9 L���s*@��N�{�nu���
� '�|�{庄��%�Rp��Ӝ�o迼K��҉����N���AkFn�թg�KZߙ�Y��g�C�q���P�2�1�q*	7 u��<V���{O�A>����j�M�,&j���xseD�h��;^h����D�Р{X>E�Yht+V��^NT��\��c�������g�w�Y���#�$�/ߢ��[#�5B�mk�X�Xb�v�Q�d���
��+h$~�S����D�B�DIٴ�ܵ>�]8��
9YK��:��mx���R�U�~w��_w�e�`��Y��J���R�֬��}��\e:����>�R���n(��g��d;��mN�*,w��~��3�>���.-��1���kei��������`�Bœ+�'��)W�+'��˧_�iu��^��.�=Ւ�r�� y�ܯ64U�t���ԡݝv��ŴQFbPX��������,0�D�Tq����?&���d
�<��)=&&�Ol��1z�MG[ʺ��y�$jV� y�:����)ts� +��u�9-}�g���\zЉ�?�j�Iv��|1M�$qJ��o��rB�.jw�_�"�-�\�{�\hr�ҝ��	��lP�:�~f�9����3��a�����c*��l^Y3������_ ��m�jk��&�Ub�������KV�7����v�����DS�jD݂ӳ̘b�#���q{/Ӓ)��(��7m�����+e^��y��3�QeK��m���a5��e`<Q�b�h[�E��<�`]B�{Ϻߏ�֩�}z�b������f�Qׁ��v�&"��!JE���b`#���g�25Ql���X~��W�s9�;	J5_7~�s�u�H�z�a������Q��8�"�:�\���E�?�� ���9����7�H���*8j����_��\"�X�������T{�|rw8� ��
s����'-y%�/6OȹLp C ��Ν.���39��0
	����.nJ���~�b����KҀ�U���=�]	{�K�\�^7׹ߙEA�U^��9f�iEx��E���&W��������/��U�]�@mdvBS&
:[����)xgQx�-J�΄~��w1ir�Xu󃍕Zb���X�釕�4  ��8�6x���{�`��i���3m�4��8��9�a�ܙ [a^����S~�sp6g�������G��Vh2�wȡ���1Y<�N �lNŽ�$g�]+���2�f5c�4u>٠�v�{Bh����{�a�?V�9:��$����!�F�����-�ڽl��b�a�.w[)^�I��}~V�ು�%�M��!�q�Pɐ�)b�ɉtg�h�i��?��N!���� .�b�@V��ў[�Ǖ���gۦv��f�4>	��c�����|�	-��C�8"a%}W� |ڥD��D�3(CE�3��g����I�=�Tk7V��^ 4�[��{�u���/��%�Yd�KlG5W�%��ŵ��?5nz�r�e�+q�B�	�o]uCA�0R�JA1ʜo��^<�m�R8�KhE���T�zdl�5X��tm�1�l����g��=�G[����l�)�1�/�856�$���*�$��u��z��e�i2T��Ӌ�<���B�$�)��X5|�x�B�Yw�ߘ��:��ekLV&8��K�Q�f]62���1n�������Y�K��L����1$��}�Zxt�eV	����� /��ݽ��6o�ş��ׂH@j�wI\0��8aLҹ�I��o$^����Q��u�����#�+ژ&.���)J����$��L��v;:E� ��TZ�&�zF bò����p;�n(�Q	c�G���gM���a^L�V%������	�O�P�Ƥ�%�^Ocn] �)=p�d�!�e^�`��%]y����6K��A�_��A�#�1^#R����P������: �l�i+�g��KVL|$k�[�ٷ|f�K��K΄��m/^6��H~�$�}z�j��M�B#�H�z�������vX��s����1�uk��O|��ƽ�s�GAbT�2?/�:,H�w�ҧXn3�@�(��۝��"�9:�/Z#� I� ePk��ө~��.Rd����B�0x3
9������2�����J��|�Gu�W^ʂ�ɘ�������k�iJ+���d2J�?�@���.Y�P�9rpc�W�%�{��Vs�{8�눘/�N�lGJ�TU�S���i?��|ȏ>=\�?���$�8�Zj�Ѐ��	�=�\j�����^d?E�w%��##}l8�MX���s����4�! E�@kϡ��*�����{ ��޴~LĻ�D��A{,s[��l!d[h/p�6m_肌���l�j#e�/��_�y�3���؂ZঙA`ф��R�T��F|�P]�^eU�k~A�o�kS�)�i���j�Ho��ߓk@�V���yX�#Q��I��r��J��KDy
�Ȍ���#���g��I�3�y�7��g��Vf��S8���Ւ?-GP���7XH㋱�zl���m��I7C��P!!g��t6
+� ͣ�&/�/i0kD����"�K�����3���l�~WM�l����v�"�`�5�55y�y���#�[N6.�0��6�t�|��e5��2��,W�@�X���`�$I�$P���	�	g��������!'�~Wôlv�[����ԃ��W���ޘoGR���q�<���fҪ�z?v�9�)Z��Y+�G`�'y�+ � p<u�nb�e
[��7�C5�.�eH�_��@c.�'f	q2!K��L��H"��&�-�G�<���W����J�\+� t��u�ꅣx�Fa�x�V�V��W�c��~�Q˫�K����!h}��?_��9KK�"cWt��S���4���CA_z��|9�[�����[����_ecs�`�f�oHǘ��#�����A��5[q.������ӄދ��,���S鍉�m��x{
���/>�ػ=��ຳ�bl�����8��]d���I����������	��:��G_fQ`�~y��-����9J@��~��&�7U�ͻ�lW�/�s#���L�5|A���3���[�#�Cu�.�#����N�i����� �=H�s��!�U���Բ��h9�#9Y(����w砆�~,?�Q̰������=4#�/�{Hv���Yy^���$$���h�MC��6P�Gc���CW�e��9T�M��z	&���j��I!��GT���v�:O�G��*d�m���b2��иX(���i�庀�b��"�ԁ25��K)o�P�tBx�מvW
�=�5��m ���� yϾ��+m�Emm�& �h� D��H�x"�s�6R�]�����q"�;�	h�̫rؓ#vA���l����ne�@uB����C&N�· o<�ш�gq���%w8M(�:��o��*olCT�P�v��찵o�r������NE;W���Yw�o������͜�H��t/����*0[�J4��o׿E^��*���p�pyv�4"X��G������^����f5wm�o���@BL����,�yل�2\<��A������a,�VKJ�o�l��.���$T.�>"�W2$&y��J��	��)�[2r�W��I
����;)�{�}Ԁ�j���i��� �%݂O����_#4��`�4F��D.
�B�n݈�晥��~�͏e��ΌOU_z�w�]�D�m��]@�ܚ�����0()ј��[5���S٘�=z����e��=�(���<�u��8<J���nJ���{|b���~�f�!QG~�2@#��{��U6�����_�S�GL�xp�_x��R��$�V��x��À��@
��I�E��`zT�x�����~�BU�8}� ���
PdAR��7N��I[�t�!Yk�>�r��{�~�2� ����E�T��r��h�h��<i�T`/���,���Tu�Y��'��K���wh�A[�*�>=���=�F|Q��!����ޓ�V	��帨q���2�K�k�H����K��R����xK�QAW�!AF���K�;%�
��7��T*�R�L�''�?x���7�fx�`1@HG�©I��d�}���2���^Wͦظ�mF��*v]�W3ȟt�Nr��� rГ�HA JqGX0j5�.s�o�3zE�XL��q�P����Y��U���yV�OQ�e�t�%�a�M}mk������i���a��Ж���Z�l��}J�M�)�͐�"�ǢP�equ��=pyb��]nVE��f�Б&%g�枎e�z�?���\u8� Xqu$2�kl]������Ѳ�T���g���t��� �f{h�,�iT3e!*����+�G�˾���y��۫���>l�{
��p�j�m�ß����!J�L5s p����c����Z��L<}�m/d7��Kiw�i+�zϖ�l� ��Lj��6�k	��0�i���]ᘽ��(H��Ur�u��j��֩�f�o5+Ǽh4E���Z��16�x�m�u�!����m.�+'���(v�� ����hp��`Ԭz�k/� �1���b�l�`�D���pM�}R�=��ӱդ-_u>��P$�[�ݪ�����;x�Y�����I���������� M/��q�CU_; ���7��}L���jp�{�P|�I`�$���0�!�5��ך7Bt3�&��Aƻ"x