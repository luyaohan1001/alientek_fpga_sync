��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��^:�P�o|�	�[���߸Y^�u�t�C��]�QCLlw"��<[g7��f5�dCjƂ���k�����w:��4�K���\�KZ� K���� �����`��uJB�� %z�#vy1 ��QC�:��ݳ�i�`Ҵ�|�&IШ�P�������P�d��S�^�@����#e��rY|�@u��ir��Z��.�HX��w��*18Põ+���U���K��4ԛئ�P���,�8zu�m��W�|��'�˵�U�2�v���1��Z�L���7`v.��a�b��.�_x�����6`�[��k����vc¯g��!4m���V��+|m(1�w�����h�S0m�T�w�t�_w���l��!�sIN�[n��jG�����٨O�C�a��Є�.�{� ����r����(�x��s�OW����}Vs#�P��o��a8�S�����oOϔE�����9%�����	�Wˬ��:γ{Γ��
«9��1+0ą��
x��d�uD����Z���j��kρ��o��	���$B��k�y>�-�~4��UJ�h�+D[�Ι ����HN@��_#�e�pU���Eԥ�V(���T�w#Ao�dɘ�h��a4T_G��~&�$ai�(�f�j��Y�n�gI?a3�����a������X��sAD��C�n�hi��z�0��	qzk��w!�V��q��o���6�=�V���? &���K!xŨ/�plؔ4�	'�g�duZ"��C�ᰨ��a
t7i���XBl`-n
E����8�u@���Dd���	��rNFH ���c�E>�2�� &����h@f��]����G<Y=����C5}�mR}!�����g2ZF�������u�Y�1����5[¾�s'9-��%Ld���PRۗ2 'Jm��x=�	��f��աJk���C���_H�'0τ�D(7��#$�xN'��r�	�5�]�>3������??E_��tQ1�v����Ihh����\���M�T�����}1�?`��buv$���=T��j�(��h�Z�LP���0n��#���>�Ҫ��y����_�����N�3Q���Zzg'����^�"�åM*�M(l�6`�R�P(�$4��h��uH蘬*ef-�b? �Hs���Y�Jq��e՚�\�[w؜�U�4�J��g�zK�VS�x@_(&��bx����AH�2X$ /�A���3�[<
�-b�:���ܶ�����Ȯy����0��o�Se� usx
�@�3*';��Q�Q���(	�{�M̦�Ƣ�[e�J4����軕R�#�0;�����o��R��L�.�˳��5><��:H���D�p2LQT����e��cUe����m��'��u�;��gL�"�V��<I[���U��y�]�x�8�����#0"6A���~('�M�M��L�Q�M*�_bK��k���Co����,-�E��h�2�1�EB�'g�3W�xg��tv4@aQ�Q��aO^�/�p���re����l�0�³(���z��b|��xP\���g34�7�K8÷�Ƶ(9*%���]�Dv:/U�W/^5�3��1%�TW>��V��B�;׸�p�U�s�o[�=���G�/�׉a��D}�ד���U骑v���;p�Յ�\#U�ED��~���5.&�/��H�Y(s��x3�q��3Em� �z�Rl�9.�=�B�ɠEkv&Sa��4_u�F�B���h���p��N���.*Q��Nܐ�_��lw�g?�z�ye���[���^7P�Z�d�k���v�O2e���s��i��l�1�R�������,r���9:'3B:gD�eB���|zq��5c4� �����k�����V�QKa\A��R�,{��#��(�����`@',��"��qJ�50�G?;+^�\�!w
q��z����}���Y�,�Q���>��S�}�;��G/s@K���̬�	u�Zߺ���Ug�?*�6\������`�Qc�� ���Zb��J%*wU����N����.��.���!�@����D��$� a){�d���ܣ��ߓ�	c �z�?Ԥֺ8}��W�H�jW�FxH��o����h�\��%�t+gYg��3St�;Z�Ę�q�u��,&����	�����cY���;��/� yc�V�M3���Ɖm�����ؐ؞E	3ޏ���Z 8�z���o�.��z#����d���# fL����@rP.q-�4��	_�5,�{�M�yi�����D��OAJ�V��u���Q���G����eRUH�*Z���;���S2~�{Z�WA�����R�p��Z3�7>�4=B6�E�H`��!�����#S��QP��PK4�!؁�����
)Ug�7㭘,>��&�&�٘I�w߇��*�%�o:�GWk�$VeU�r'����KCkDkL^���u
� 2� �Pp���E�'�*����#����������{��x&�K_�43���E\��ALf�";��5*�g���kw�l�]�m��#4g��Sz|{]M?�J乱�D�1�ډ­W���'j-��jx�U��'�����@Kn���Hy>ʛuV�{Ĉ����#��y�;��zp7 �vP�cO�%���Z��,�
�z�>r����>y�fp/��B�(�\:׼���~3�"RH���H�C/��s{VK����� ��Vi�F?�rE�Hge�}��-Y L�`py4���sDq���A]{43i��YDY[�$.rb�6*��-�^����qW{���s�j�a`���y�ͭ|�2X�l�>q6��N����*Jw6ġχ�:�:zS��6��#�Oi����v�:!ݖ���&#{zg?t kf�2l�j�w�i.��)[�>O�.��}�ϮVeQ�������v�c.�b5�{3�����H)�:zLDDE��KR2�?Y�rt�J2)a��gٖ�o4�۞k ��g%�_#c��R��!�F`o�zރ��Ƣ�Ő�K�5���M��W(�-hO�8�NA��e!8���rf���5$� �E�0�{�NJ�._��Y2�$6a#�������ۘ��\���l	�)Ͷ�hu�I��UԚ��A���x���"�G����ڜ���s�w�#	��fB(#}��>g�{PQsi��~21�:��	�mw�s�?���*ӘĄQ���?��0+�|�k�(���j����;|#|'KP���G*a.������f�l'%j��<#ʒ �p"<g* 2:�׏rk�����#��x��B��� .@C�I/r#&���_Tf�ST/7n^b��s�!�Ȫ_���ږ�ֳV4� �(:>y\� �h�q�%#��{���͆�K�\��zmy+�d,䥛����b��*1|�m�v�L>��G�%Hȇ8���v�w�}��c���{1H��.�7��b�*[���1�V��up�fg�� m
���[r-��|���])B�G�����o�Q�&�74ǺYu��1dtר��{��y ����!�«iǑK51x_��D��@p;���ƙ�3yg����)��\>�]7����hGZq�}f^�D'�Nj����ӟ�t�p,3�v�)��ꯑAk��?V���Ȕ�x\Mg��A�Lx���u���0YW�2�a�B  .��Ϥu��K"ON�lT�S3�����h����I4=`;�!��NSU}��������w��2�4Ma`��
`�V^H�m���D��r��w +�kW]Xen��Dgɇ�����1J��K<��+;g��S
=ZLSn��aTK*���8��U�Vʨ���dRb	���
dTٕNҼ[���
�fa���b�\"��Dⷺi�ΌɆb�䤑&��̚_��t<#�;���cSe �o���&R_M���`ݮHP�x"��D�I����g��A�,�w��s��׿��$?�b���������f�K�yõR��ě�����_2#��M��.�/�>oܥ���6�Rp��Y�9�n�}��:}Ԃ��|	������^�1�v��1Җ���\��>7F=�T0��, su΅c�H�n�1>`��7D(��WË��0-��,ߑ	��o4
ZI��W��/�h.���˙x����~+�'�"�b������j�D~
�#��x�x{Q�0i0���ѯ��"�ϓY`���ME�,R��U�d)PӚ���hAY�Lk�9�hWg���{a=4��>��� =2{���R�7IK���7;5���쵓���z���Aa64;�PC]?�v9�{N5ϻ=����� �t��t��v�ҫ?�q���Op*�!�=��{��L���F�,�ej���;���,�fP�}_nZ����\eP�:;!Q��1ݍ\��|�/�9�K�k;�A�������Y����I_���ԗ3���`k�0Q�J�%�¹�d˒������w2*����v?��p2��֐����+�ڧ��g~����φ`��s6�mđ�
�	y?=ߺ�����+�h�"�F3 G���	,q�s��p��M೒�t��MYE.����Ֆ$_}�:Za��;�pA<-�D�*w���J6����Y�Ҋi���#t�7$� �_�����7gQC�X���N�>�Go���5/L'n?I����.j��4	x�3�gM���y�m<%��0�ƋU���}��ʿT<i�����ۦ���z"���y������Ϋ濓*�X[Ns��x�I% ؾce��A$Г��ԦH?�vD��{��,Q=$�¢y��s�B.~';.ֲ�k�zk�먬A�ݴg�Q��z�Z۔;݆J�߮Ĵ1��ʆ��܋޸b�燪��!�2Ҩ����[
�����6ӫY��}anSCo����F��o��"*�`�O�%Tw"��Mj�+�� Qy�f��;˗���4���<Y�`7��@&��iy�������X���!0o��HT��x��q��s9:1WKe��fx`��h��ć���A��!u|x�\$*��~�Z��0�uBy��Q, J���W$BD;O�ׁO�dJX����q���0|�x�2V�X�3].�~[b0=�;��a�s{���,�<���9�@>I9��=E�9^0%�"<g�3�*T�[�Q�~�� �����=wrMg��
�,���"���(P�ɦ)�L�tɦ��wĹ����d�P}l9��=~�A�\�[m��
�?~I�v�@4�5Rr��p�����}�G>���N(�_����l^p���q܆���;i(�0+�Ӆ����2���\;�kZ*zׇ�+���ְ�e+;b��ŶlR��$��b��/���x�V����x6�G'���v ~&�*���矤�4�AJU�gYm���f�E��C�;�lg�)����wD2I���]G�4���VHxĝ�:ݔIB�,����wh�`� m�t�t�����,/	����L%}���m�������N�R�`��<G��!��_�t�̉x���X��L�3�4zލ�����RޑE��g�]e
��d�n��@���ZG)���`#FJ$;��E<��,�!&-ۓ�������(wˁ��C����T���Æ�T`XCD�u�X��^m�j�Qv(�={��CiYT���O?��L�%��$���F2�%}J�b8L�IN�]����_P٬#�-T�9T���^�@R�>Y^���S��8�/���./����IKӭ��n��ڀ(������g����uumXA.ne[T��!���Ԝ��n�χ�|�����~���A��1���ϩ��)S�o���G�Ճ�L���4Y�7�S<q05�	��E�p��"7���T��մFe�h.�>�qy�������������kV+�B��@�=��+��h�x���h�0���T��i��,<r*d3��߽c��ة	�U�l?�_HMg>����>X^�/!�'���J&��Y�� �|�� ����������5"��̟�=�|�v%į�ͮ?��<Fr����1��lXǌ]*@,��}ϭ���b�U~0��r���_�5�H��EZHW�H�}���t�\�~�{.(�JV�wN��l�I�f�~�s<�%I&*��;�n0���
U��{�M9�����o��x�5��ET�|�DM��z������{o,c9,�M��a�F�b��+��Sq������wS�e��Xݺ!��'�6T���Nԋ�SJ���.ɭz�{h��������}�����v)mb����C�*��J�-Ϸ[E�P ��������M�y̟p����R���t�$!���H��;���1�!ȑvo"������(���hf����|�"�B�$�'߈[1q`vO��@��*zX�m��]��WEt+�h���C�����Ĝ�,���`�Hrn����^��>��>��P�W[L�tp>X�_���;;��/�?ն�=,�r��(6�X���\�Zf����y�/�b5��ϐ|�)_����=���) d��'͹ƚ+�6^��ؐ���jf"�e��/��i�����/����{6d/��Q�n^��F�R�HtoW��7,^���wS(�
�{��P�%<K�緎������^j��y�<��M>�T������o>�EX�aޫ�e's�94~�ɞ#�!C1]�d�=_?������L3��M����^��S"��/���%L�Z5mfw� ������h%���#��@����,y�K�S�T�MuM���Yp#��9	n���P�u	��͗FR��+��:K��q:���Z�4x��7J� �8u6�	b%�wֲ}��^����hᨾ,�m3�֝���Y0�*|��P�EW;���םkS^0��i"��֪ǲ���<��~[�v@`3��,v��8W��	��J�����7|�Ѡ}\5��%��x�@1yUx1�-h+"	��hT�'���b����Ho�vm�T��2�mpI���	�Y����"�\�z�
�ѾȃZ�R�DQK6��D��ꄲ��Mpm��g�:>�3��EDv��|.`�K�9���!���7H�|��_f�iU��1�@j���#�E�{Ot2����eSl�TxhV� ����ФĢ'�,��q#M��&�����21�ncy�RҨb&	����J��oa��ZwI�Č���|ԗ~���k�l�S��F��|�10�4��(����	�A���$-??n2�Ϧ^Ig���f�z6�zh��Q������b�0Э���ئ�]�y����.����U�Vr-q�봧	���ЏT綍��xTU����y�o�ӝNod����{ro4�v�oE�U(��V^��Ĳ'�������>B݅�&
�+k~mI#暑kk���CF��WRTK3��Mv���X݋��<D9g����;;����*��Yp3� �	���I���8xi2�+��˶� L�6*��H���m�Ge_=P�K��8�[��(��[�^`Ł����4��tvS��Y��յy|���<6n�`E�_�n�S�)��� ��y7x�� ���x�V;m	�0Ҩ�47�;W<�*ׯb��; QԯtTX�����0�Y�� l�,���(W�0L�dp��DF�S	a��S�+�	�m�����Ißzg!1�Uy3Pu��R�]��TUcL�$�76!���8��qE1zֈ����7��2T�����˄��a��g�����l�k?7(��M���0͢����E2TN����FeI[NX]���w[$�W"� �D{���}7�G��ٯ�H�K�tF#�p��6\7->L2�
992�l��P�7��^�G~�h�u.r���w���Z�݈%hX���;������o���@%ƍ�w.����WJg0�i�Z����w:��f�TgV���.�(WR���	@x$5:���
�m�(���ڡ� �����ǌ.<0{X�0mVf�c�|`�e�1{�k[+g�C�MJ��xB~�j~�ǭ�r���wA� �ݿ��[�<Wl�4y�f��s,�8h3ٻ���	Q֖������ؠ��dj�`�� DnD���Ŭ�sč�v���d�V��qkD��
��k�I/Qɘ�h�i�����49�9�$ |�	��5 �qa�RJ�I/{h��R�����x��{0R�_r�}�(�Q�ɘ�G�U��	]�@���3��)s������gP׃�	.���cA�T�""k�[���tյs�5i�=�6��^f�u��gH�X�����k��}V�*�@K�ع�YQhb�9��b�z�`v�	�iMϚ}��tps���Ѫ��E�+����_��`%m�dՂk9��)u���ֵ� �����=#
7��.��phA��R��c#Us�>R�'��O~E�
76HR� ��w���lM�wwj�y9��WF��kf�"tzryy�]�BxOB@Y|Jh/3���� ^I�҈�5�4����d�V34��/�Z��}�Bշ@
����r�$��ol�A�qb�_�`rY<�,:�K�� �'I�	�tA�K��/<˦}�%�p}{��=7���K�H*sISbO�G�BE�p��X�\�QcWh"�4�������9
��u���b��v�<��0V�/3Y�w[��db;�Q=��n����,���h�V:���hn�"�N1������t*�ȭ>X��\%rN�%�XbY�gCB"��so�'���!�u�'���f�p��b&��ub��7�M~l��mK�'5��z��_��=��z�5T��MB6q�o=ı[�[W��.�vrp`�`j�	p}�*b4�����'ǿ��ʗaPw�m����<DJ���ȼ:CZu����&��X#Z��LK��R�o����nˉ�|݂/�A�i�#�ݼ,+-�AݜТ����G5�'ӛWyU)�?-�eX�\���b|��:�W��+%� ���h�r0�޷�Lq�F�yQ}�L�"m4���K��b����?���G)o�فQ�[x��>I�r\���T���U�_�e��	y����]�{N0��D͒	',>����E����[p�p�' ���y��tY���U�Qjug<h	tI/�q�'����������5�x��*��7-/��/(Sb�8�����l��r�`k7��Eԏ�`ZLl{�p�Ȳ�y�xo��8Fw��(�#��P��	�Y�H�c�^�]�z�9\�� �s�V��#yG2�|�X)w��ki龷�)�\=5�����؇Y�+�����]��_o���e{����u9��`��p�>�%i�f�;ó����&��>�� 㓍W ���ZP)c��	Lu2����\(1�T.�=�p�:�N:�����ޛ��Z�}o�+d���u��ƍ�X/ʯ�g���TYBL%�8��~;n��@�F��	\�����`�эڢ~���'��߶Ao��r�zu\+���qN�����.j�ߛ�5�����	�k���J��S�٨�BJ�ZD�Zے@D �{+�/�v ���P��a�txИ�~y��u9d$"}��d���WР�7����js[�1rX yͺ�v�ٹ8��P���Bo��xӞ�Ǚ�[<�>� 안dcI��ȱ�>�)rӶy T��L��iwG|d?1:�ec�!`�}��!p �����T/���Qqx�}�3�)!�$�'
\��Kf�i1@aW�3�s��ܖ�i�z��Ǒ"�C��S�6��/���h�),�ǡ
6�$F��0A����֚1��d >��A��)�R�#b��T	��ȭW�V�tK���,70��޼��Y@_���:�vMW�_�^����8�QCkC����~f�~���gx�>��K����_�(�,�n�M%L�7����4zay����Y�q�-Kx�a���$TJ" ��8�{����\�q7��c��l]R�^�jc��P
��o<\� q�Z�G����9g�,�k������.�vQ�����,W�š�`q�(� 5-�'(vd�fs��tP��HM���D㓃�.?%{$�2��,ۋ_�mF+}DW��T�?�ݸN+�*T!��h֒�[$�+9��d��%�j�#^��V���Q����P�9թ.ZN#M�@�(Ey
и
Ƶ�5�|�e��sa�wgy��՘乪��ؒ��0I��b���8$L[ȅz��8���pՋ�DɁ4R�z1ߥ&2ϼlu��3o����_������j�w��N�"h10|��WA�o5j�[�o9Ayx�l��D�9�`����c�b�J�I {>�Q�qJ�gm��5�/`��
���$*�Cq��vG���<��]��Vzq�m}�[/�Ep=_����ݼ��j�K���NkKS��剾��z��Q_\f���>e�'��;��v��]}wit�m�Y��	�0?�"���*7�5Ǻ_�W�w�E�v��
C�g�4z�5�~l�	���n��CF����@�4i�W����/e�j�Œ��zo���y5�hzw�9�a��I�MϕPJ'-0�s����NfPGf~���.��43�nY�r]pGH���n�6�2�=-7���4Ue��n���ؤ�U ��_4��\|�6so���k�z+��.j�A�yD�*��~��~?��BAE+\C�[53%:�Is���:~�mj�1��9�8��mwn��&�ʹ����&h0諼��������r�S�&I�$!��+V �U𙳔��G�m��|�=�ϼ��/�T/G����-^�Ϛ�,�(]ݗ��bv\g���1;�v��H����·�����d@�5J'���>' -��ϼ�a�ÍNX��1��������w$��S9,�h�ܴu�i�k>����<���$����~���R�[Da�C=e��8׽�N��Tъ�x��+�Xy<����T};��v"�gۑO���5=�Ҷ8*Cԉ࣌�w������&G�DM,_�٤-��8����R��+ǔ�����H���r���K�Fv���������I�X���)�@E��n�'g�-�3��xr�,A-d+��r�u�XO��R��b��m/����{�6�$EV��Ýs7
v˧��%��M�aI4��/B��oT�O5%��}
�\� ��$P��ǐ+t0&"�VU�{.�C��̗��q�7������`'M`C����=[[��3�A��z�B��nZ߳L2w�q�ȸ� �ǰr�_l�J��-��(��������1��\4$ �q��IU�'J�;���W�/z���Dƿ~-mC���Jh�g	�g�o������8�[^��Gɐ-re�01��y�ӎ	��>��,��  �5�6�]I��@�m\C(��q�(繈XeB�no���]k�{_���eN�m%�H�C�&�e�rJ��XF�t'��k�b>$L\�E�.! րe�uBi��c��w����_Ѕ]�B ����G�-��d1��I�O�N�^+k�.�[J�ř��v,�0���,� #%�2Da%�n�*�_��vs5�2%"��*C��Ѽn��[�%Y@U��*f�=L��X>�}"ⷌ��P|灚��yͫ����l���_]���'��o�R�N���E��RzQ�uL���: �h��aB���1��>!(;������ݶP<6h�'ࡿz|���'�6�g����8��ɛ��T�r���_�4vE��3UY.��k�b�،6���?�~����Tw���G� ��IT����	|"��C������`"\��_:L8�D�l����O} x�[���]��_�kK]W��kD=��(����2ŹlQ����-��B�Fz��S.�q�S�S�m�`�+��g6�����*A�4��ҧ3��^��F2�i?��)����%�7Ok����H��������Lb�}Ӫ!���㐪�kuZbm�1v��J�ubBXR�G���B�*�d]�t��o8����av\_ ��&g)��=����f�)r�T�e�NÄ�5���vn�Gwc�<�{�$�mG��0��:�ג/&�ꝇ�zk$����G��C<�A���H���{���0���t2�w�2|Ǆ��w9x��`~�"��82>�?�w�/���]�N}�9���]��dQJ%Ǐowy�!|�A$�ϥ����Y���3P����� ��N=�(��Fi��$g�n���HK�����MrT1QY�0o$�I�}��WQ�f�Fi(�z6��H ��	'1ۨ-&��/M�Ӏ~��t�6�S,�L�_�[?�'�����|�B�SʱJ���k�7۪(�=��3�)t�ivDj]�{u�Fg�"��*��-�q���Ǘ�I�%�][�����vx�ܔ��Ͻ���4�W2�i%
r]]^��	�z�|W��)������X��<g��g0�~իbY�! �!rN�-/���,�oec�̅�Zc��֣ܬ����EC-oA�ANDOR�-M���|Pn:�JF�8�(�?K���A'���UXZ,R���/	*pGn���0���l��_b�;�ǿ�E�P���7I;`\���E���?���ʌw�x�,���3�y�����a��'��S�Uc���+v�	�����Qe3���I<] ��Ȟ�3�a��D���1��8|C�*�ߒ���q"�y�<��c�M�Az�3�C2@�bJގ�AwV�ugJ��-q_�R���'����U���>2�Q(�D����D�%�P��G�)Ϛ|�K����{�z�7x��þY���hj)��$.���	�b�B�oy^,��S�0"pHo^���xG��2�ڑ�[4�����|�ʒ?��m�h� � %��7Mm\"�I~��.��xE2^k��6)��9�[�࿪*~wSC�yt�5�§�C3���bl��'�)��$�O�U9�]�>h1�ch�ԡ���5�%�� DF�?�^΄�KbMy��g���!ّ�rz��k{3�C9Gp3�kߌ�i��mJ���D>�7���B��R�ҽad�R����M��)�s�ڕ}F�$�����P��s��y������p,ꁂq�*��]��j�N`u�KX]b��Cy�/��#�U�����J]:ϔN���b���{]'+��J�7�H��f���ޔ��q�G/�g["��.\���tN�v��_���'Z�����7!b��Խv	,zo�/�]W��IQ���h�O�u�Uz�]	d?O�)�� >	lZ#05�q���оr�\/�r���+r$%���ɫt++�?��}5J��m	���p�'��!�<�L��۷�5�A�<�
	��(�j���]�J2�J�x�l�g�'�b/�M�1��{����O�ki�-���*�(�D�^��/p�:���S��k���55/�&��v���OW�V�ҩ�ǒ;3dآ����w<�rr��-qeXl���L������`b���C_ӟ,��?G�2���<��WXI_�N�e��hT]��o&�e��1j� sA�^#��ѕ�MN��2jM;~�l9t�� \��������K�R��+H��zr��@���,���;n�yB\W�IAA��fUP`��a,�I!�W��n3�ӟ	�3v��rZ	�_I��)l�vkw$�1ͱ��r=�y��(� �xѠP��L�/<f4W!���@���0�ud X2�Mׇi������J�� ��?&����7�ʼ�u��=�{��ߚze"�٦G�R>x�o ���"���G)��BW��O�<�L�<�юW"f!n�R��&o��?������~�&�Թ�04H�'o}�y/BCH��e�g�JZ��Ewz��F����Zvo�37*�u��	�<Ur�eCX�(V��q�~���)��U@��&��٨΋1���u����bx�d5�����]s��^r;�cy�xЛ}��!�Ȼi��W�.z��]b{��v�5�.���idC��g��߯����+q�����B3Q�-�Oш��3��<ń� Xw?���� ��>:,��ׂ?̠%Ff~_[4KN�G�e���Qw���]S%c�;�me�}z�k�E@:��D�l��\��GZ�+�)0&z��~�$���:;س]C�e=�����l��+L|DJ��h��8y��{�W*�������
���@N�!G��_�8�T]�'��z'1ո=3�Ә��Fd˯�~�υJ�����^���;��9�v��[P��z��+o�(���U6�ȧ�ߐ��.��n�:ԣ(����%v��74;��
*^�L�2h���a��XV,4���ΡQp�o����AcD*K�D�B�
'�WԵ�]EⰛ�S��f�04ϲ��:�r�Uc/�b�V��|�y�%�7�F�4fޱ*Gd� f��}5�7�r�P�I+��*5�E��D����Ђ��0����K��}�Ċ2Y���4
>�r�j��1��Q�>�ܷ�����o7�Iߑ�R�8��$T�1 �]�.��kNGz+�@���H� ������}u|H�1��;�����e�A���zK�^2D�ch �4�J���������3��Hj ��]ښ�/Z����A� ��DS}3'��Af�d[��g\1�u�nz��s��&hs��*s����-䟽��;?L���\(�����9�P��a��K�P��^'�l]�}�o�^���#K���Xr{~���R����]#8���xw4�;������S���=�V�O��w��7�H^���=|�-w����<�6.��i�,��T��{�6��A��t*��0���V��
7U(�۾ą&뇈�l1��7m>$�#�=�c_Ȟ���
#�3�R�x� l{�-���ݟ��騾w�RX�TԠ!�*��D�L���5������cv���g�3�t�^E$G,�{}�o�ϑ�Ŕ���7{m����2QgA~U��Pm�fIh�'{
��+}*|���U��`r5zd:�
����$��;��gs��7�<\�~�:N�-f��hplX�A��jQO��lQ��9��~�=��)��-1�?:Qδ@������H�V���i�X����k67�MTw3�U��
�-���wnw�ژ�#՗ţ`�!�t�&����#��)��kE��:�':|�M��JI$4�ZG���r��h�[)U�$������W���AI�Wj�?��H�Ǽ�j������6�a�	O���OP�=�h*O���o�Ԙ'{�oj[�zp_j}s}��}a< `��N&���'�%n�4��eJ(H�o?��M���(��L¥Gh����>>Ӱ
"bx��p���5��`|�-"  x�'��!�a�-����W�����]���F��J��O�(4_o���|�7�٨��	?�n��(���X[XF��SW�f�=h��E��w�aba�+�=P�'�r0��B��>M+?�|��)�P�<b�1�B>�g�CL�Z�<��~�N�%��}|;�/�߮��ޜ�Ҷ�,Z釢W@w�F�8��T$s7[ ��g���ǘ��Ki�V�&�bXq	.?*��W�粳� �n�fR�(���~�r���'����[��N]�V`r�ټB������կ��M<m��y�0�����b���x=HEz�%}K&@�:�����[O�R��?]�1�q��-qr���@��L2-a�eL9���"l��Wg5Z��,�1���F4S�H��(�Pr��W�T��KH�m�� 8��SS���et�lp�b�"�b���o�^�����_�36�r�6x�����&5d��dY?;X�|�y��n�96�a��y-C��ŭ-��{��8Ā�9���OL�5VS��-$9��@�l���x���	vH]x�r�Q�"̳��v�ynQ'�%=*X��ԗ=�.y�w3N�)N�`��=R�^]�;W�D�V��$�[�N%�P����UL�j\�2s����)�Q炉���'5@�������7Ub���q�Mem��8
�"c����⒅�������6�<o}8F"���]\WcY<)3�QJ�]���2���������Ԃ���i ��@9X;�z�a��Z8�Ś	ȴ*`�E�Q�����|��|�S���slm�R��;o@so����Xp����7j��������ru"��3_@3PǽH��_�`�S� ~���o5k�.A!$PgW_�����;�͞�n=��n"�gš�}X����W�^�?+|��+M	�[�Ԧt��/�W��A�L�΍%S4���v ��c{eʱ���^�*D+�R�Mg|�����P
P��y���ͮ����q����lF�̰*p����#	�X�_�5�!�祣�����e�ߎA��U�ɦ:�m&7Ye��#�75�T(�("��u���<�M�D1��M F�ʂ����о7�B��u��)�I��g&_G����S��jp���h���QzcER}xe�x��nJ@Z�s��$j�I������V2�����YbK�yj0�-�-nwNi�L�9J�pY��5+��
��Ӡ�/��B�N�1��֋�[U��K����Ι�x�(.qO�q�������y2�H�v�A �ϙ摠���3��cp���W|5��<@6y�u�x��sgqj8Ơo�h��m��հ� �\����c'��w�y%��)9�w�Bĺ�n�kv��QF��vMy!}֝u��U�8�Pn�Ol�C�r�4�F�[��P�
�B��s��g���� !Ac��%�=a侯u��L�-�B3��Xh�,��FC�&��w�X��V��,�4upP#'�O�Kme��+;��#phӇAٸO�3<����<�Ƴ:��]�S ���/%�X�=m��_�=�<�J�ڞ�K�21�r���h4��v��������b* �o���bȤ�Qf�G*��	9c����${�/�`�`!���>��Q�T8E����z�����\/��|j^2�x�e�\x}��jo �����ڗ�&��XB4H���.�ݍ�q }���q0B�m*���e%��ׂO����i�1v�
.�42�5j�Ҋ=N��ץ�uBx��Z6���LV�:�P��a�B#�F��]Z��/,� �>��î|�.���1u�ս��9��Z�틛��j��5g�F�w��au�H[�!��_�r�q��7r_nҡ8�)|����F�p�,覟�t[�YS��Rk��K�$jhc�Ķ�F�h`z;3�u�}�%l�۫�^E����\.黻��Y NE>�X��f����jɕ���p��9�Y%5�K+L�GΓ����ֻY��(M�'�h�͆���4|n��ڙД:�r�)�_p�7�U��E�Ɇ��;��-� �<����r��m�ZՉ��Q��Z�=���K
 R�Q�/K��(�1:$�@?{��a�|xTƱ/�0F6�˹��֤O��x#��+��z��-�*�yقp������vE ��	���vg�����%v:�Lt������^�:����^���Pk������]R�}j��/P�DN�a₈$��>o��b���+�-����&:�WݙaP�D[��e���se<��8tu}Nr��<�1*X�~�Yx���x-���m�Ȣɿ"}j���2|ȶ�U�	-�פ�����Y���j�Z���=vVs��XOkc[�jm(�8!��8	%*_
�Hs�3ؘ_�xF�n�kj��E�w@�%%�ªLZ��p�A=�}pdHO�!iG��3v5�|��r��s���e�za,�x���Z���_` WE��F���#�����uI.V������M��u��!��΢I~^��
�ps3^@�^8��U�ǁ��dokA#�(��nz���æ��yG�&H��t*�����B��_�d�O�oː��@�p.�6(�)�`��Q���̏�YZ�& ��������S�������m�`k7�I�ݜ�`%��(�9vXwI���݆�)4���ٔ��F�ZN])� �|�E�T��o��-	����-��*yu��rѥ��)Շ�(ڨ���s���kZr�բ$y�3�ބ�?L垞4�'<�c1�����׵=�7M��yѩ
��߷���u���݌fft����AF�8�K��f�N���d�I��16m�HV����#�Z~g1�ף�ˬM=BXS6�(?��n}�'?�>�b����ɑ$Mp�u�/e��9b���X���=�p�:-mt�ψ���#�L��Ǧ�X���1�^�\bǞ����.0��٦��Od?�_PvY��3���nO��3փ4�LCU7���`w8O��n�md+�v�vo�(9��n!�Pp�8���lHe��} �����=.e���?�T��6��p��f7�������Rr	ǫ3��B�Z�1R�z�Tל��M ��[?u��
Rэ�{��K�e��>~I��|Ijf@{�3����+�
�S^�C���QtK,?`��e��'O�N+�o��gX�K�ά��J�����S�:�|2�q4v@?1z��#�'���*!����HQ8��e�yd�8~9�	z�;L��`r*�ⶼJ���Y"<}��Se�zt�iی2��v]�Qb�y�X�7��ví��9��J����x���W��`��;2S��<���N~�)MM"?����q��5�L��	���D9�IX]HU~�)%��Wz���co��M\�tT�w�I.��Y*ފO^<���@F�ƨ�Y�GH�e�+���Ƃ����%��4��g��g��"SB6����,Z��E`O�8ٱ2�ˎA��?��=�"�=�e�yܜq�1X���8M�4r�
�2Q��g,T�sW���ǰP���&�{�j�Ǿ-�P��op�=�d��@ZF��+�+�8%��-_��9�Eĺ��|&l��>v$D"{gVh/��&���óv��3�\�x�gE�52ED��K+"�9%�gU�89�NjP��)A���Mxp�85;�1&�'�$�K!�	(L96���eW�{1ﯮ7P��\�9���A@�.�bN�RsY��Sg��{�^+g)��i"̃��M�'rv�ԜP#]7�)`y�
�{�w�P5���Ɍ������^�#V��(���0B�%�,TpmO����X��_G��&�#� }�gwTr��p)�oL��u�*�0f��ؒ����<��&3��0q����]����iй�1� �t���/���.Eb�7�����T�߀��!�{L����'��<�5|/���M���[��WC�[fR�A�xCZs����¡�jX�*�S����<C���<V�j8��6JN�sE��JK��H�2�s�F��ڡ���6��U,~֧i�sAqI�N��X�(�h����8~���+���N�ϚAu�HVl׳�k!�arLhE�j\T1�:qd�o�U��҇h| "��;Fe3�������3:-��+t�@�M�:Ԍ8?f�L���~M(�Zɇ��a������&cG���BVO��"�*3��X��v��F���H�{�D�`���r:�C��X�3Q�(�WGc�"����a���/��H�ٰ�ͦ��7�'��R��1���~�*Mc�ZS�=�t��I��y1�h���?Y�*��v��(%5j�{���m@7��5�e ����Ƣ��"晐t�K�u7�	���j�G���q2��h�&!���q��J��k�n��Eu��g���Q�Fүz��&-����M2Cw�.�mj��������x������x^��m�5� �?�`�	T�]J)���_��J��*��G�U��d=�c�Kw> ��81�A�ҷr��R0��(ܗF��Q����x�T��Q�5u�yر��m��#_wJ��A��)�N�Y����3�\�-?â9�X��Y88-C�h:�̺ ��_U�� ���%�wF2��+Q������S������v�,u�C]#A��68� e�
3�w�Ą#"��q�u\� �R���!B���Z�v�3�	J��V��n�~hUZ�!�D2� ���u2�,����$!���]PU#���p�0x���/�:��v���G���.���-fW^:}����k���'�ʿ���i��ݽ:�I�7#���o�iN�q�(
RL~�$ڍ^�/����S��D[Z]%�
w�C���`�:�}�~4�*!�[�������2})SX!�H-�Dg��%���˕��9HZ�RK���J�y��==�y����8H�q\_.(dط�܂t�'��<�~�_)�V��~���z�V���]����#�u_O4'te�޽��r���h�6�c�����\�������)��σ���A &Z�7�l����(��@@↛��Cr�K#"��#������V/�C0"�iEe�n����%�*� �}3�An���c���c������ʐ�#�.\��Xyx`3��uưe�E�7�r$ z��W�R%Qԙ��cwl����b�JL��Ռ�ʏw�e@pOc��N����R�X��ڇR�b����_
��Z3�`���)L.��v����>���2�Euռ{q���=oEص��q<9GI���_���p������_5����[�
��$�\e����6�п�[���B]u��b&ho�=K6�ص�I�(�(}���ݹ����lh�B��6��<oq�}X�1u\��B�1�èNui�uѳh�VI���l�15�3�kEA� x�踩T1ѐh�.�.nq|����ש����
q��kp`�F<uk�#�h��x���a���7P)-���};bi���\�'t��8��� �iC+Ʀo�t��Xv\X�kN�0��'��9c�����p�����r���US�P�����W�n��8��sU��>��,�45�:)r�u	?���nK�(��h��HJ�Xbl�q��,�Ǆ�l�?�~���㤉9h�[>,�� 簺ȼb��Os��Ex�ԇa�Ep;�`)`��,�7��0�!��5PI�4���8��������e��m5Dⓙx�y�A�� �@-X�ߦ
��?��H	dc�7Ū'�4꟰3ʻ�~��&������+(�+k�/�E���3�'�zʿi�;��yaَÛ�T6M�%͛hx$a�|6+u���`l:4�ʔ�엎��X@��� P�MZ�@�����j�Ѭ�^S��P��^S���ſ��O�K�b4���:��5eWa!�04v���d���7>�Ci��'�#��U��+�7�3�|Bn�A����m�u��m�1Y6�+����s���KQ��
�Ir8"�4h�i�@����%�ؽof�r����e���|�U�?�T(�+�����Q�ߖ-KVP� ��.F�r��ɿ�J��p+?2�	u�q�����sI�Sh�ߩ~�E�����[�ޮ�s9���P���4 SȪiYɉ��� ���FI�� ��t�"�}���O����ȳ*&H�3���vH�3�߃���P���Pu�A�4k��Dnz��2�i�F�q;�ɺ�[�l�8>����y�6�J�9Ʒ(2hG��}�N&q꜇���.|#�/�2s����R�/'�ʣ�n�)�NC� �i�:W�]�#��__�������{:�X�މ��q�z�WJ򸳽��2��@���e�A���( �	
C�3�TL�(=�����Mg`�
F_�׫�%�p�X����E�{QHfX�?,��yi��Vo�P}����4f��eG!:� �n��{n�?��WZ���iV[�O/���v�`j�o���dn��gX�?�ӵE��b���xY1��z�a���%g�{��bڽ"��@}ۯ%�ԉ�Z蜚]�����8�Pv�s�c	��^�<Qh�ޮ[��Q�*{�y�PF�pM��-g +k?��|�T�GȻT�l�)��Jg�U�ԠR�����~�aB���J�� s%z��z]5���d�y9������X$���Ô/V����MC5��;Ŏ��M��b�A5�k��t7n,)�b���(FH�h^��������w=�(5M+߱������o�N��R�B ��ʽ�g�w�o,$I�ad�%l�w0���b3�ޅ��q��T�R�z�O��T9�*}��u��i�|�.,�c!c�\��WU�#@T�{
;���H��z-����A(�xaHt�����,�a��&��QG�v���X��_ɍ�A�P)�W�]����j�������5��O��G&)c�"�*i#�=v���8��`y��K�����%�^)̚��@��XU��+���E����v� 
u�:?�`5�i��9H<W]3�YZ�SÙߺ�5�hb	��p~ ���TJ#�H�a��03����vRd���-��5����t	0��rsI��"l� ���BK�C�������7�e'6 �B c�)�(��+�;h�V�>���K�[�䁡f���p�@�����lP; �6Yma�9ZL�B_�|~�?����ga|�b�[F���y�fO���4��&���B�(�q'�tu�ܰ����e0m[$��lܛ��3wҸD��ּw����v&O���9i}Tе&�O �4���H�p���k�Ѐ�Fj�
1�-ל�@���1�S��*J�y#_Y��K��V��jƴ���]Lo5����(��b�n@�bw܉#�/��b|E4���LsF���	^p
�������G�}Kq�q� �+�$I�.UH�7�ދ4�X
i��s�`Q���/��HbV��A��»�1��h�iHP����W��6=�J�_��|A��Q�لd�`��ȫO�=�Mc��o�(p�W+��G�䄲��7o���WȾ����6U-�W�s��ó5�g��M.a�'}������(�TsnV9]�t�W�9��@���$Y�Tb��� *�&��Z�fFV	��)l�����E�MR.��(�����R0@�xڬ5\�u�t��o8<�}�-�@�k��a7::��پj2�	�B7����zN�w���1�^���p���M۷;ȴOS�~��-���]($)x�&���͕Ǽ�&�U9M�[\��BZ��t������bb�ZޤCH/��6�i_���j�����RN�#$�@?{c�HQ@4���n�&J ��IZR�F�S*̖1\�/�1\#g1�<���tM|+��v�K�XV}�E�&�����6�5X ��k��<K���<$��������V�en(�lA���M����q+Ɇ�[z���@���
d�K�8���vc-o�;n�+��_l|�1����@���F��8�����*UH'�E��#-ȘZ<._i���g.�x�{�:���]!��򘀫�C�k����hDIBT����N0���z��K`V��s*D�����q�17��w�� ����z�J�C}�Z«?�U�y߫Dc���cR��sliQ�hR���#&UbN+�HK��N�yw���UJԨ����i��m�7��5�WҬ�5�Sd&�To�@qE�˻�;�i�.�E30�c��APW2�;���V�{��=0$pI<֨������`	��4�w1��ة;���a����?{J�%?���k��8�l�հ{��t�|��l.�WGìBe�(��U�	/ѧ�҄�5�e�l�n3&�	�|l�UV�lo��z`�f2k"j�p�~��[�<G-�ޭ[�5�A��(���c?c��	r�y#=�Ov'�o�&�X^�����B�]_�٘���qD+b�c����F#�E�)���lݭ��sH).r�N}�s|�!��/�w7���3� ��U��ф��g(g�2�� Q�	�gA�_��"��#D���66[.� {Hr�� ���ne�q>v���,�������aF`|�j��~�i��B-�$К� v��q�&�冏z���D�#�����W����?Rn�!�&�nɤ�>�*�u&`��<*��J����v���ON\��e�y?)��c�ye�Fr��|4 ������ܪ�'6ܐ��o���M�@:����Y��Z����;d��"0kQ�a�;�q�g�}Mp�О���11cS��/��1:Y�[��K���K��[F<�����#�Tryg���[@ޅ/_Vn|��S'��2$�4����~��^5Y6S����N�В�pkBq̫m��~21�@�1ֻR�\Z����(Dr����Y?�(��/ˌ-��#�K�S�Ei����(C�~N���dQ�r��HJ��V����������u�]�g`}��g �pX/�d�ױn�����9Ʉ{z��j+����Ix�Ԥ���m/�|�����A�:��X=vN�ݸ?̶��Rcd�}�׃.��T�n6�<��i��!�U������|��7��-$}�����Q�>ai�2e��|h�҄Q��%��=�\]�F8po�\���|����).bm��8���<�������xN���ы�qb��>�I�o	9��W�gX��$m
�P��b���.�4�l�%Ӣ��]���AH�:aډ��U����rrqK��e|�y�hjw?����h�̄��~�G~"��Q����P�3��f��q �
P����q7���n�nb�u��w��6&���(EB!���(����;Q�`�$G���`�ZI�w�bu��*n��{�p�'B{�����qX$#.e�g4�G#pM`�L������Ti��SFʿ��$ wԶV�\�w��|�������2*x@:���$�u�x��>�>o�Y;2e�+_@���!��͆� ���f�k�U꥞7�����)�J�C]M�1èb�¿�5ٙ��.a2~0å<��QQa�}�4����Ro�$1a�<�Pţ|����p�\5:�u;��Lʓ��@��%�ӽ=٦�J�)++n�#Vk�RQhT�VJ2.�
���	@#/��݆�lBE�S�	����=x��(�Z|�r�T�_%k��u懖#g#X3s��}��XQ�"'���]�	Az@tP��,���?�	LM衾sK3��e�D���K�z8�]�2�܏"� ���PMA���8!G8N����ַ�g[���.�`n?�B����҄;���.|>0�CB�^�f��^��{`(bg�Ms7@�Rf�0�ݩ���,ÿ�慖o�ʜ�~޳!�v�P	B������)H�=��q����(�C�{��x|�2�#��+iJ6�p�격�C��е҅\^\���h��ک�1Nπ�=|z�7�%C�[�--���b��� �l�%��';z��Ȑ�B�K�~�^ k�dSyטQ��}�'hʼq���H9��jWg���'N=�m!S��^�Zo�|�#&�wND�q���:�5]lr���F*�ACg��َ�"�s����?C�G�k�R�PÄM�k$�[��<,�;��t�Rh�ٌF#�k-S �R�2
TD�RN�3ac�<f	���<%q��G�:PS�4V��[v��Ag���*��}�ν��Bq[;U�-N>��k��t���tR�1���q�T�soП$+W�΋H)7u5��``���>��׊��p�Ϟ[:87bÍm����#\�D�n�~Km����D���ʂ���BD��8%��\B��2|��#�|��	�e"�cFMKk.DǗV�ꟲ7a���"<�SB��%��{-�Ǳ�9+E�R",� 	�J1o���5.ǣ2�|GIU�\��zH"�M�=�eHf�+���J&D��5%~M0Qk�0N&`Q�RDo^�Z�B���s���[R&���S�?�W<�����Q�Do9��Rc�[���z�q�P�t��)&��`�,�q���F��b�R�x���q��jU�5�g:�ˬ��.���qy\cȀ��9�����Ѥ�i��9H�&D�Y����#Ӷ6.�>p����d~Z)�Z�4x�vO��+�j�/룳L�:�@���O:��ΎM&��V�\�p�Y�r���M�_t���o'd���w��6�'��`��?R����h���ҽ8��9�D��߹N?��''��=�|�w�3.x*��R�xKS���5�U,��ȿK�r��:ӀVlV�ـ����'g�ՈK�L1��}0Hח�5�Y����`��>3�,xp�D0�e��Lͭ.Y���wWV�Q�z��v[�����Ǹ0�RI���`����'�b����@タ4P�Y��~�5v�-n��$��Fr*������%�
���s��)4 ��w���\��8Y�|��3�0 K�)@ڇFy��R�i����:!�g܈`�����Y<��+*�є��SM4���j��\!��& ��O���G�#,�ʾ���>�ȑ�9�`z�x�eud}�ᨓԘ�J��qN�a�f^i�X#	*�$�yDH�b�I��񂵋S����NM؍z��,�ޢ4�B�h�4∪����#�?z��a�Z�eޱ���U����r�7W~�ӥ��� i���¤o}h^��"�DH�(�I^�`��q�|��/�?
\U�!c���!gޏg�Y���5�;Bg>�v��S{D;�rW��!��N���_#��B[DN�45��Ch��B�J�3��@�I�{
�Y=l�u����>-&���T��V�$4�g��3�?ꮒ"�l��%�>:��� �L�r�E�qA�3{8��)�<�\�6�L ��PXGD��E�o�	�"�������"�������[����3t�ތ�
���(�,��DNף���j� �^��L���J:ˏz��Iw ��M�Anw�n�nMM7���ou��5�(0����2c��AV�/�����o�5�!Q�ZxW�o��J���������i�����\�ۖ�I���l�e
}͌���@�D���*|@�ݨ��P��R/a��e��E8Y�s~�� z{�/{C�D���s�N)ڤ����eg�c��e�F��LYn���A���(o����߉P�üT�U8E�Y���Wn��T�sr�Ag���4TD�ʋ$���W�ڤ��7����:�8�ޕ�S�����AHyy�]k�?���x�[(���\5I���xj�KN9BA�o����=�'�mI)����m��zY ��}9��m�Eo��8>�򄕂[��@^�8��Ɨv�ͷ'#60��$��L�o8�A�qC���=K�fQm���K�9ʡ�a�iyWS�VL4����6�}d�j���ij��,T���]Ś� ���u����l4���AK����ƕ�䉓Lo8F�`n��.�j�����d�k�qx�[���O9I��s�9�4����F�����:�.
�ʊ��v*�J�A�K��?g�i~��tV����S�?"Q�]�(��ŞzJ������#	!�e�Y�R��)F{�9�gY=g��1���K���7V�j��(ోk��E��T�%������=��=}f�B�+�+�p�7��,�|���.�5*�â���[�cN�����!.��X�[���q���Z3��ʄEb�hQa_�s�L�4÷UZ�WFj���6ħ�?�P@�?%�Cn�E��S �Iߙ�T!��&��ݓ����-N��/�3h[YPst-�bq�w��w��rK� M�Z�*of��r�yw���G�o�B� 8]�	'@7d��9]�� '�"0�p��Ǝ�_.�Ai���L0'Яt8�@���m;��w���T(}H8�5����_�)��'�<6tߒ'w@GV��Qȿ�Q��V����h�?����p���>"�u��S����LZ�7L�t0Ҡ�ݚ�t��OIg!��~rs�c�x��а=p6��C*֑~߉����ަ/$�q���8�N^�;�>�����p��r#[�82� �r��ݟ:��VCs���|,�j��c�2�>�7p��H�F)=4�1<�[EK��%��ͭ�74:Xtem&m��߷�JM�P)��e}K��͏9������+*�m�If>�L�cV|����\^�� b����0ܒA5H�]!���z�uύ����|����\q���B����E|���Z�P|�����óʑ�C�n�D/�v��Rf�o8�v���S����p�ƚH����gYD���Oyx��,�l#��j>]y�^>�c�#���ԟ�]1��R�'/E�:Z�P����	���`ڌ�_��S�"t�Gc�"t���	*�����6����"�����4Y���r�>�y���*>�0MR~cl���$���6�j�k�����G�+�v?n��F"���=yI���:��$�8�w��@b�����<�m
[��c�q�r�7�\.24k�Ȗ3���v�k���:��)���g���h���2�	_;���Cq�*�3�by�/*|�
�"�%��I��ޔx��t*Y�
�Hr5������B����VF�^���d誣�U,#��hTuSA��Hr���(v~߷���I5p|�7�E�,��0[��*̤���0(N8g+߳`�)@Ҵ� ��PQK�Σ��p��y�c� D]�X��g-;v�Nf��hgH*�"0a�P4��J�ٮ�t21_Q���\P�ȣ�A[;�GgJ��L������h���t��R���J]�f��:_ōy4H���K��P,��|%g��������i@�t�ZBSg�U�^/HE{��֘k:Jμ���)��0J���z-g��ˇ�I(�{(J�z�3����H��d.[�j���*��if/�@��Č�le���/M_�5�c�T��{�yx�߳��#���;��4o��]�eL�N���U�C��dm����a�#%�ĀXK7�����a������3m��HpAduƈ��CR �;�Չ������ܗ�if0�5{^�i����M8��h��zb�Ë�~�K�����p�2�]=�U<�i��N���6�`�_�K3�
H������;H��:�:}:�&޻B������,�Ywn��H܋�]��
%�f�S��D02"��}W=ݓ	s�j 8�����I�M�<��|�T꒘a�I�V�ڥ8���FOP��?�hu���k��	�Z*ܾ ��a��o���X��܆K�V`��m:�~ߦC�+`]8��p�9��i�fR+�ʥ=y0�>+���F��7t����d�)9����ފ�r�.|M?�-�侠�{g���g�>Lb�t�?U�U�E��U|1�)��BL�\&� \N��*�~Swe�//O����Wf�6�N|�`&�m~8�M[B�e`��mw�ӑ��OP�������_wa���B?u*�B�Y"�R�l�h�1����o�/�#X���6$g����TVu��vW$U�)��ż��n�H�TL���3j�cD� q��(�)��͒���04��I̊�
D�S"��_/Z��_
(Љ��s��|��������#��m��8���Ui�>.,0�	�S��3t��3���U܋�^J�w߼�*����?:?�)<B��<���f�eS���%i��K��6v�Oɚ�9�m�r�}z$
2��z���$[b��KD��$�ب���i\9l2��N�$��%+�߆T�����J��4�NI:f6缥��+������gl�u�� � &�^�C֑ B��7;|����a#�D�^z���;}�'yn�s7��<#��� čU>�������,��]dQ"����)��W��'��g��Nxt��M�eы�-�pЌvSج����&�'��瘼��d����p�*}[��R��
�zuE�<�z�*�qbs��1��R�Ij�B�&:g2�W������PJ��V=��dk5��T�w�₾�P�v�����%qx�)�	�gՅ���}
�u�}
�����/ m]g�M+<��1a�oar��C�t�`}\ݑ��a!����F�ɬs�o��-9Qz�s|��a��9�PR���D��� ]�%dF���Y2/x��(
iT�[�%�c�N?�v�VO�W:=CH#�#�ܦV�[�tɼR�z�����fm���Q{�$�m���m%���?SA�,F�)�\�5�R���D-((1���ܔ�;x�'�B<���F����H0������3̟x8�{{���,g��$9��/.����
��/LS�P�q۴�"���q3����\���#{�ԭ��m�"��$I������G{s��I�;�k>T�O?������$R%%���8%�`���M�����7"�{�8��g���O��dk������\8Eb=ӕw�'x�?"���gi�N��E��*�%�͍uVq�Z}��[F�Gb&�>[��*��m��g�M��\��d4.[�� Z��LmfS*�f*��r��Ō��e(��[L��3�D]�9���4r1f�>�$�B%"��61�s{���/��8WT,��d��^�K;Wh�F����"]�3ᦄ�^ȷ(8I�%��������O,�.�7�O�� bHk��\�kh=�8>3���<'��<1�v;���-���>}i��l��C3#�:�W��m8���v��j�!q�F;D�;�hyJ;��m���
�x�oc�=eEǟ�MOy�[�r�/�z젩�'0�$�k�p7��J��IÆ�� Z[欉�}�� Ÿ���-��0����L0�y��`�z��,f��Nsg���p�v���t^o-��9٪h�G>�}��N���N%L���*MRk"�j`J��Xq6L�>v��L�$��7+w~���S	�e�FWIV�:�&�N�JX΄��_�;
h`3j����2������F5*��p������!9�^������}�hoV�Ʈ��,�Y�9�g��#��Hs�k��SҗP/�t��E�ZQ�-�1\R�P��-�� ��������1�M�b��ۻ#�U��!�g��:�N�OC���<���w��^XʧŠ��ax���zI媠5�,$E!�?s�>ϤR���Ï�$8����&��b�'�,��0o��&�4��ɶ�m�T�-BdP�u��N�˽����jk��׮._!(N�G�ID�w�|EF�h���SP*`���j!����ǥm0Mt�D����q;J�՚��-뭐o���T�^DD%E(����8��v_�.��u��ʇ���������`��?��O���Dx�����������bO�;������.�i�U�`���1�!���ĥŢ����Ƿ�3�E���LO��x�b;�>�O_��(��sn8@i�����<���#�%(�+�_+��׻VRu" �n�Jì��^RO��Tgu)����!��I�Np�u���\ڃ��)n���/�D�3�N����WR��7������E
�53v���7_0�no��C�E^�����\r57-;.>^ͳbk]��O��d�z��c:�]�vhَ2�[���
��
���Pt�]�����1�`�yP�
`D���1�C��9��t�[��臼q:�W��}�Ξ]��g'4����Ma:|�:ϩ!ť�=�2o��5wF�d`�����5:�J������O.̽xͰ�}��C$`��Y��m���ZN���9}j��`�?��HQ��JTu�uZ�Um�2���l\��8�v�j�آ��g�.��Z@�ӳ�\��tA�jCsA��
E��ь��~�����\hv�Ӵ��J�p�����]�����f�ys�b��~_�������2�	��&Ϝn$k���_���u��d;z4
ڵ�A�C<�%:�;30�ٵ��22��g����I��u�d���'_]4��Q����zs��n���lϮ���0zQ������w��u���m}B"#�+�d�nԡ�zJM��#�8�xWa""�#t�V̄ϒ5�@���,O�>96�	:�)TC��iZxq�����c`�?LP��?��5uqL4�z��V��6Vy�b�ٕ��Y�Q���v~��W�t�� b��i2/b�;��%�vnCoM�G���T=���_ �,Ve!���&@9S�F|F=^Ny,�O�7	[�9]+�����A�q87�`4[J��(Nz�"���4+3�r~�I�n�.O�Z�aV�����Z��K��m�y��}�%^l1�}xhi�}��eg�㷸o�c��u]e���(l)����b�~0�s��0vJ� ����u�`�xIXK���9_Q#�0R��q�6y�b06�k����T�T1��;e_;CaO�]��Q�J�
��n�V�i�w�U�8bO��~Ľ�E^��Hqн��S:�(�Jdd���93."�-���ٺ��5���y�(Oq�Ϩ��g����`�j��dttu�*�H|���{�b����R��p	p3��6�[��F�ݓ�Ԓo�л�w�	��^��#v������2���+y����7Ny��yr+`´)-B�D�ﱹ(n�-��a\����ܓ�j����߫;.&uU� um4�2���U�c_Y��X�d�١~�8:a��������Өi�!%�C6-l�6�q�BǠ3�A��f2��{i�y��%���A��XĞ��X���B��9̕{Hz4\9�.e��N��w�SȢ��R��]I����BLh�N=nF®�W��֮1niI��ER-����3��߇�U�:��R�y-8Yhթe�^R6��oyŦz�2i�6�?��*��n8k�P>�|��r�[1fg�íۘ�܍�#��k�n,/���4
���"j��7�<�*eN+Y�|��lP���x�M<G��e��V~��V=]6�AZ�ؠ���9�iIh���:��֫�8h/��iܠ��g���������u��n5�j�T�m~������Q�d9��v	��i�/�R��YvZ����0}D�|gZ�8\�F�KB#i�
�_��q���;ZF:�S!�Oѥl��eJ�h�z	��D<�T)�վV�C?+����l��dK��:D?	���a��j�qx�Kg)������{7�<o\�!K���=���$|�\�~���؉�wu?n@鬴����"�����`~�ԅ����4�qb�5x��A�ym���<�_s���vjp*��j'�I,d>.�K�jJ_H����?��v{J˭S�$�Y6��(�Ћ��'`@��D�RD�F|��_ҝ2�N�H�3����M3�X �}�@CN��[�U2w�� w�oF������"�6���e�b+�/Tc�o0�Xp��J�8�?{������B"=Xv�Ӗ<07;��=k^�܁%�3�$�L����r��f�+�Q��1D��Iv�\���w�1����s�p`{��R��R,��P���Y^a�C�)`��@n����ٶ��|E����FG����rF�&~i�`Ǿ� "=f���~���V�3�E_��12?��ȍ����2UE�5�֯C�[%���L��L	h+���^d����ȞU��R�=�֕�t.׎����%��]V�cȃ�C�.T��MI�SZ�%�l4�٩0ru��O�(�j�>t�4:�{�0_�gM�/*	�֢�B�����b�aLavF�P1J\���|L�����2�pև�(	�t ��:P�Y�̍P%�$Z��s���]/ڛf��]9<��_�[l̑U��,�$�Xs�#��T{��,cZIC?��%��w��4�F���/rߙ��oz@����w`�wM�1�w��Tl�@����j���b�Z���cT����g������0��
	X[A�Bˋ���#ۻ���N/2lQM�HvhG �E(��s�{�A�Sq�M�zZ_��:vzS�������#��勒?E�2[PZ�7�@�[L{��Z=�B��i6�\l��Ū�RU�S�k�%�\r3�1,X����fa�Q��q�(�s!t5�Z���ʹ��d�{��>U�55Trܢb�>l%�	�P���?�E6,�@efT+n�<{F��ؗ�8F'G��~����BU��R�yQW�?�$1٬�?O:��bZ��1�!M7��w�S���ʾ��y�����p]{˪@����CXkן�v�T�����^+�G� �Ux�h���սz�3L��=��"L�fgub�^(���O6C��Ai
1���=c*�r�*m]	=b'm�t~v{A�яu�c�E>jA1�SE,Ļq��9W�H�iFb I7,�T=�]홑����K{�������=��)x���,a	/hc�=I���k����?͍�-&w�$L�NO��h�
���Mg��Dr<f�� �I�S"8G�~��E���iþ>�@(~5W��	L]��<���c�?���&{�5�A+�������<���j��q�J-�&�o��}0`%҂�:2<�d�X�������4�ZH1����48RI�A��ʲ�H�$K��>,"�F��L��'�0Vq�9��tB��0���<'/��eu�N*�5T�"`�Fp�-B)�4G��.�R�'�Em@v��E¢��?!`�wV���#�;o��e3�Yx����(��Pь��lt	����  �
��h��G+i��z�`�m	�~Ky��P�F�J^I��~nLX �1�k�I��;��G�ìKnWg����iz�qP�rG�Kud<�x-Ƶ"m�@Є9���t%j�@�qJi���Y��cfa�&����"wȜ��R}��#zϠ_{"\3�)����Rg�
�Mna-�(�z����W-��Omg��;��&�L��ӽW���I���4�=LH�TI!{�2Q��GY�<7
�N{��<��ڼ����K�����u⹥[d&�fR���{�����h?	hJ�2&�|�?���tV	��&|&:m�Av�k��A3��# �C]'��kK#KІ���A?޾Rt���T���K��Wqq���!L]�v�)G~q�<�@C�&I�_V�b'Lw9xrb#Uvtq7y�$	�c�k�^`�+�.�D�l�h$CqH���d@��Ug��T$������qK�qq�<E�|d�4�*��~�T%��ׯ����ž?�P�y������n�$�^yyŵ2�l[����v�(�Uـ��/�������o��߀���f��G�wF2
��q��Ug}'�as�+���"O�kZ�¥\Q7:��$I��O#�Md+^��T�ދ���:�Ǵ�=����Cv��~ "�~bߨ�����Jן@��A����7�<"uF)�zԎ�(l�� �vM-�ȓ�Q.�<w���:2����� ���9��K�V��Л+�bب#�D��������'�DA擜|p�Pg�I{M��Zw�{<�;q7]��O^���ig�_��rr<���ei�N�g��ٲ��<��/e]shhT�kh���CP�T�C���(0�tfzϢ��l���]�������l�{c�yx����EM�Ys?a�5)t>������1�́����!��:-����i�����]�|�b]��V��8�F\�.�:��9<����t~�pz�:[;�[kM(h�TW�d6��$O:|V��Rǩ�[7�������̕�xu0d��	p�)y&
X��X��p�]w��5��te�rY!��ڴ5�d���`�L�*f:UN��G��
�������w��x�1e�Y���k��p^��=k
��|V׮aMOg�j�bm���gZ��q���K��ir�#�{�3���	�~[_�p)_0�8�+:��k72:9����z^D��ྡ��K��,���񿴺m;;�	����/T'. ����:�F����I9=�G),txu��L�:�����ä�-��!Y�e;��k�T)�0ޟ�$L�k�>�kF�
�/K�v�ģ6]���Z� �=�r��Y���. H�R�Cڙ0�PqR�\	&�?�Gt�4W�|N�����ia�NQ4B���+�k�KU�����u�.,F�M�C����K�k����v̽��h�`1�9���eT��M)ioF��������EG���=����A��C���
�=���O����^D1BwN���_�8�����Yo,�Y�^!6�� �,���*���ƲV�l4��@�j�uf�2�����eg<�:���n��3s����?j�{-��ؙ�EiZ+�#�o		v �>`n4�Z(�ח=�8A�����}�c&.j�ip�5MJ��������H� ��1���[��_u�-�6vX�-Kz@x�E/�]$ϣ�=1�Y{t?wH�ƲA����2)Io�z����@�P�o���i��p)]bnW�`])���mY}:Bl���H�̑s�H�^�/�~�)O�tZ���|me�JwI��EO�ڂ\�M�g���EIA�����BX
��=v8������ՙ�F�X�73�z+\M���H�o4��.��H�#qp���.����e�N�i��+��O�Ȅ}�w�6����Ldf(��+b4�F��o� MÉl�ʕw���g��\tMP�����P ��{>'_�����:+��Z�����c�ii��5̔}+���^���0$RD�\3ֹ'�J��u+�o��5W�})���\km�o\-���L�A	'/�L��aOUZ�f!e�0=֥�ðt�R�pیA�����K�k�R�������)��צ�\�-�k�{��؂=���з+_��e�E������EK��]ƕߧ߁���ށ6.\�7�@�<l���W\�ǋ���o#tZy�Ih����/����h�4S�+��5?}��X�M}c�MMf#-i'TvX��0�z}��ؓ�t��=���Ъ����/�T��/���3��=�������W��(*�	��u�jsB�]*��~�a848�r9'��$ItqQlu��*���x�����$uU��Asr̀�B���,[�&cLb+�j����H��� �h�����.���S�4{�2�;a�kLS�"�F�!' ���A�34��*��Ĥ6x�I�;�����$�O�.��z��+(�Yx�`2��J�LZ�If�\��]ѵ����K�YX�����赽ճ��p�������=ӡ�o9�k�L�jq{-u��bWr�J���C����Q,=x�ϳH)�r�X˨@	��	�L�\��z�$�"1*�D����4�a��Jv=��&�S`���4��vtFU�)��ū���d�ك��fE��5�Ȱ��F��d��M��~����/���5=�L(=3%G#�1{�.���ukA���|𰭼���_�����l�v���9�(�����������d֐�J����|V���-����L��TN�12^�Pa��J�eK��3�b鑽;�7O�٬N	���<;�F�su�8�b�������Ț����mM��]u�G�<T 7p����r=h�;�ee�.I�%�`"���'U�����:74o|I���غRi�!�_3�q�T�\eS(و$��{'��+�#x�:{`�x���x���S-��V���	�A���ǤU�n��S���VR��b�b���'9#7$��\��������D%�\H��]��[@Em�cG��;�Ѹ��R�\������'���� �h:G]M�M��	e0��Թ��N ��^9�����8�
�d���/�Wȗ��ɻ�T/�o=���DM����j���Y�h(�s�5�β}��
�6.�6�.Q�/bFF�W�hϽ�?�g���54Is_C���ƣO�ˬ�� ���	����nn]�jE˧�0�Yѣ;�'�}�f���]%�E	�7��2y��(�<��逴�\����g@pn/	`'+Z��G*��f��M�6�V���8�?g�#�x�"zjo2���٪
�_z�lAk@�3�U&�Z�U��pW�
��R���.Δ0]I5�A�ђ}h��#���`p�`��h퀧Ԝ�6Qa�$��4J�;�Tŏ��KS���pDVx� ЧsK`��_^�m��ZZZ�˽�Ҙw���ɽY����d�
o�ݑj��<�$��FIu��T+�˞$_�7� ����5`+n���o���r?�t˻%��e�����o�ˈ-��^��J�C!�oR@4:{^�������^^��|� ��������W҈��wB�Q���;��#vn��9T�%q+�h|n'8,�1K}��j��e�~�G�Un��vG�y�ǋ5�*A�$=�RV�%X�����[��ŷ��q�ǃ���#d��iI����+���~�ǐ��d>$�������)0{���Ǟ��ͭcC��iLpg�P�Do���_|s�<>��`�Fb��(C$�Sk�Fww��r�$�6P�$�0&]:5�h�3�UN�H���3
x���2�!���{�2���J�Жs��\|mH
�6BʈXE��m�qS��Hz9o;iQ�pj��߰;�X 8Kh���L�piB�~`32�1�Pq�ƨNPc���S����ƺ{#�+�G��ơ��Nu/��4��Ň�1h�����	@2��GA|���v�1 Ih2�0�ys*�	ˮg��1��u��e�G�jJ�Y]��C�ߞdO&��SB����w��l�;i���4�#�j�B4��OF�- �z����gٶ�#f�􊏖HO�lyh�24STw� V��t��{���K�ԩ���!�H8-
�l0�b��s���Y�\�sU�r�|�����h���B%M��tެgV1���1�{D�����[�T�_���w�!�~�e�&\H���sv�Lɼ��~v��-�.��������)�!�t��ƿF�l��ocj�30TFס��J�=?_>�����cRа��-�q�t��R�6Be�X#�����F��&ֵ-�rFk�껭u!f�O�-�<6�c��ķ����I�q��1v���0f�r�V��}��UEb�~i8rb��ރ�Qa�v��@잣�<+w���������l)Vʒj���>�&�H������ߙ����Q�����2T#�ˋ���0�u��}Z�cj�\`6e��v
���O+zK"S�S5�9��)����ڮ_�k{0�m��Je�7��/���8�p9{��\������W�F�M����B�=![���[J��Z`>Dn�M���"�����?71��tW�Ch�:8�K-�A�lc��-�v�����R��l7j�O`x�Shr�%5Rs�	5��:���_���i���|�Ӊ�|k}�^hF��I���]����`�p���[^V�zC�w�j��fD:*_�5�\`�A=�v�;�������(K���d��L��_��'��rR\�y��g`>�Au2�
&4{���Ơ	��E<Xy�:Ɲ�sb;�rBDA444^t)���2���+�ń���V��E�g��]9�~'�:�u��@J-�Xçh�+
9���2f?3*��o+`⼆��V��YC̕IMvBY�6KZO�&Tf,~\��	' dЩ�ߔg`�`�){��7=/ԮWNFa.^���u�)��2P�qm�����&��K�Li �i��������4�\a��h��-.��ϔӽd��En�L��戀��Z�C!2��o��`b`4��R��q������|�A	�8��OO�n#�h��#���j�v��t��@�Ȓ{�P4�� ���������D�z؇��ē�ŕ#2�H��T��b�V�ڼ��%Ic�N��BFvg��<��y�-��㢵S���T��J�}m?����h�¯��pU�nF�f�4Ni2�%��G�iyu _v��2�}#=|[�+��?w��*��	gHbG�ւ�9Bo�V ��h�L��F]N�s]+ �˛�EhCA$=���u~����I��ओx�d-@�;�\??���v�L�X��2�r��y)NB>@�2X�rF~.	tMr��].�Ы�l�8�C���^�ó�5[*j�k�E��6�.(C�t$�܅���N��3�ja������MQ�P��B���>W�LKw��e@<������<ڸi�yP�JKh��x�*��t�-�zK���̆Ŵ��~�!U�sߦ�-��*5�)���L�D�>�~oM�Jd��V�g�5��vnHnR�1<!�oP��|�3Y�1�xG� ��yf�JGg֮�&Bi��W��C�쀩�:�a��U�
ޑ)�Ǆ��P�̡����I'�����@z�T�XCW��
D���p��B��.\���ay�N˿��#n=��/1���mDֻ�hо�4���[
�d(�bE�h	���Owbq�?���N�P1i��i6N�~Ŝ��T�L1@�\~Um%XIpN��A?�?B�B�""3�T���tZ�){�u�4��%\-�x�f�b
q��w�DH��b�bco5�t��������ۙ��hD�:�C9�J��6I2��I�����W@@�� t�����Y)�DJ�^�o��pqJU�=���4V���b�i6��>�#ǐ���R��f�Fʪ�Z�P���0B�M��Q�IC�+J�^QWv���쿳ʙ�-c�����V���	��x�(�B�g�0diȱ�}��Նm���E�k�F�rL����m2B�Wvƻ��,ѹ��/T����78l�l����{�럻R=�=VC_�b�瓁����\��H֗Q�s�ZE���=xѭ+#0��L����Z����$gFo��DZ+�r���o���dS���)[M����\e_Ŵ�ۢ�g���n�����@�c@��s�wNGe9�޿����_=����7#(�>k���L�ut��w���U�,��W�E�A_7�ԯCƵk̜xa��?kIK���ʋ�*ҙ	��Li&�ߝ���+�]	d:��k*:-W2�����v} S7
"��U�e�Ҟ�A����ƇI����(��rʶ�yC��LC����QqO��r/q屔��:��9�@����x.-7��<��D}�@Ĩy�X��	�f�"�bT�ݗ��Fe�0��wvX���D�A�n�8���x�l/͟������ƞah��V�$����Br��=~� w���2H�+E��8Ɛ�A�SK>��n|y�J*х�'ݪ�t �WI�ND=N��ي�ۍ�&��4t{`�io�'��N��"Y��T�W��U�`���\�ՌDC�;���N�U_ثqŐ���dPyHW�2���O�.F�=HmI^�7�� c{�l�)xj`�5��������q/m���E�H;�o�t��io2k��N��
��`��.�$��i����)�L~>���c��y�f.��0��O�/� n7�`�b3�^�{�ռ4���06y��כ8��)i�6_&ܹ�����X��Z��#@����s�J=a[�?!e�.Ch�<x����c�������j|�3�?9����Vm���;J�5fT�s�_�F����7J��&��z�S�1$\j�'�l>�}�eEmU�p�m<hC�7:�9of�:+k{�J��7/w#M�|����ٕ���>�u��2hQ�6�h�蜢�s!	=pB���}JM����?�Ng-�
*/Ǜw�<�9����@���C7���))4�`��d��z������
m����3#>J�D?��U}XB(��:�RPY��S�C�ż�!y��5��[�o��^g�ov=G;�k�;��L�9	����	D�IK����(x7�R+��74z+�SA�/6��3�w�����<�;�\/H}��4��{퓭��sR"4rw�d��K5��������ۘk��ITĘv�ԺWL3�|.�F�p�[Q;��4�ޗ|�uA�76'�����7��)��; h����Ruj�dA�8@�q��s�dIU�j�}�V[��ÂV�"7}Z.]U$�f�t�r$�W��I�!Sx���C�Q�/�FAO4�����7QR�>���I�ɴD�����T`��2r@��{����_�<\8��}��K��lbh�L}�0ե��e:��!Կѹ�. ��y+J���o�M~���h�����LF鐵�����i����+��*�F|*p����3�
�S��8�T��;~�Θ���'q�%�E��e�܍�����tqL���I�8�z�^=�ol�898Z�>�����{i̷"�.������L�Q�ex�=E�G?���~|<��`Eַ'7��è�+.�_w)<��4'�9��P��1�ڣF*+��y��8M�,��"�S�Nz�R�Y��[�C� �=r�w���q{�(��c�9�y��;�b|������j��fd����tC9���Z��_h��2��[0^�Q�w��.���d�+d�؀�}����s�}�P[.�q�M?�p:��*(�gr?��c"cOpa�Їq���%�YD��.1�r,م�7	�(W�3�
~��B9D)NS���!:Hz��z�NN��0xW��_m9efR� ��>&��	���a�Uv����L�Q�]���i� ���`��S���ci^y���:01<�L7�ṞS������	�v��3 �0N�
��N���?D�I<	�g�z�O��*aK<�����,;%Ű�v>@`�d�kDm*{�p����|��:W`�g�B�IG�%��`�w�*+E�x�����Q��\-���2"Ë~{�
f)@yl���	��}���t��+�r��I��/�����x(Z^�j���>���P�&
>��6X�Ln�/8,N���ǀ���JA�ԕ��4��z���(j��縁H��6HɓJ$�F�9/�(�jW�N���͵\�.WX\�P��]�T�#��
�����d�E����j./֟U�"�kxm��*ɇ��5���͛��7X�<�?��\���H�f�N �*E�A���	MXH��H����m�O���_{6�@�P��-���'��K��{�<K�|
���}����}b	��W�����n���/�y�J��CH��g�r��{�_�})�,����!'�]v��:x)y[ i�t&�!����R��Ch:�sn�	�DŤ��ޝF5�)Sy��]�����_��}im���B���k���,1K���fn�?-âF��6S��l*R�wFuI>�k���1[I��Y�#��,�����[[|���z�7�kh�2p3������@��px��A���ɒ�0I�♎PD�n�;�L᭸/��A=���u�6��`B�ny���s-���x�A�<&%��(�8���$# 2c�"Ӫ��h�8Һ�3o���Fɞ����	E0`��(Q�Y���W���	�MNb�ި�@s�R=�q tF=q�|1�EN������}�I���Pnq
<]���o��-��{^N��c�oUn�ɡ0���Dy���J�潫4��<�< �g���fwұ�8Z.D�Y��K�\$@�~!g�}����� ���NL�Kk[5R�8�~j���6U���^s�`�@��j���J'N۔\�Žk]����iF�ќ\����}:��c@���΄�妯�{�6�S���s�H<���d��|�[a�H�����|ƯJ��m❝����g�#fh7�\�4H�%A�j�i���N�r [Sl��/X�K��)o`�ϰ�()�� �Yc�|��fV6vN�ҦR����W+�
����뺺�\�����҆�o}S�X����}�����#�f�7�ixP�U�-�d��b�',��	��s�5u��*�ց�&rl��3bk�WN�\hTBϢ2�2M�J����%r�B��;��॓�'�e�(��y��(6q9���	w�^�!���6��wB(x�]�,�k)�zP*Q6�H2�C'������^��l<�_��h1q��1	<��B���B/1�0#��V��ܾ��QLa�2�$|WR�q�L�M~z�_���#��r:��
�>O�mv%��κ�,��ݘ[bi��7_^��zh�r����� �pA$���vA���^>&�0�#|��:�vYO*K
���(��=�6
ib��C����&$����E5֙���"��	��٣?/������c�׸i��-��F���E����ʿ0>"?1�@DY���$T���n�q7�&���3�:ł�B�z�$h���'��1š2�8~^NUmt��Y���y�Lo}"af?�U>��`��y��R�o ��Ƞ#<��9�Gأ^�J/�|�Y6�r�kcC���2�u��0m��)�����
��g�%��aU��� R_i5I;��� )�"�*ԛe_�}�3���4J����!��_A��[��ܸ��T)��ۻ��!.�TkAc[��o��l�!s&�$�!�-�8��e�!�N�g������hU��Ɉ�B�����igT���v��٪6�I|Ս��C׈���7�'�I��]X��X�n��F���7�n���ay�,�|T��W������7�K�'2����#!Ԯ��V��3׸;�k1��Hz��NC ���[Ir����>�3g��Lw�Yh�MN�����r�(�Wd�)�8�������~!Q�O�21	�`O��=�i� I��}��`h�����7�)hR�~�G��f�l�G�%=�c��NQ,�d�Jd������H��r h� ^�b[i������,�%ϵ5�)��?�)��.dL�Qh�R������7T��������N��@��׃FS�}�c�'e�%]������J�hɵ-	}\Nc��<W����sC)t�k_�v1�w�ڱ'�Ak�C�D��~�{��Z��:ꊋ�{e�q5K7���$DK�X���,v��+Yb�e���� �8D��A�|�K�;�^�e0�����	��W���������&���8�ȭ��H+O�dS�:�rk�����ǢXSf����j�aS�$�S":��Ml��j�6'��(�|!�?h���7��hg`;8jF^ήC����U��~Ҫ,Φ �d�y3ΊO��I"l��u0:S�Ф����7��f��}XS���������'���#
$ڑ��{H.��?���8>tǬ �&Ɋ{p2�d���gHdZ\{�R��2�)��y~]�{���(;�'#2L~kw��,��W��R�M�M������-0)���p�#�&:g��%�g���]�_~��Rư�v�M[p̪(�^�%'H�"���!,F&���E�FyK*]��%��J���H���9Ң��L��#���م@�7E���/��\�Ja1��?��6�aޥ���R���#L8C��$���_ԩ6�z�EU�:,���:Ɂ���`�R��ֆW�r�J�)k��)�R;2��r�}_vߕ�'���_�����( À�� �����0A=��IYą��8�wP�͔�$��-� �OӰq p�U;�N���߂����K�Ai-��*W�Wr�� K.��P��������.�J81hB�Eq}xY���(ػe�?Y_R���r��B�Cz<�2H} �+K�>��d���q���A)� Sꏎ��0���.R��6	�BVwJk�g�3tk��mƃq�B�v��zy�xY�w�h�K�S�����N?�06Ӏ�R��*��Bj�:���$mo�٦Ƃ ���.��I��q�;I˵�XV�~���2]
b��4[������}2t|�@�"f#��P�m������B���~�"��O0;$�gg�Y���q-�����Qy�Z2j����<�$�!+֌�} D.xJ�	Ⱦ�'V�1��� 3�_���|�əo(��7h��B���B�ٔo_�e(�h��H��_���vȞ�^��x@�x͛�a�OI�b�@��<��M���2�c.���CϜ���o�*%��^J��q���2hǣ�A�{zZf�H ��ꖊ��э���Dn�Ȱ:��̀k ]���_��.��&�~��}#��V�M�G_'ț�$c�_y1*�z��P�-���$[s��pG�{hIV��ll��xDN5S�V�A0~�x�&���h����M���;Ҽx���^J��;*� �U&�������gz���y!3 �1ԆX�.F2�P�W�o�}��r�#���8f̮���-y�,<�b%:��/7��'�f�<<h���$�t`����y"3���6M?����xU�So��GE<Z� �#��W��Q��Sb�����̵��㽗yT+�����dq6B���'���޾y�?�QT�t��+��0����w��ղ-n�Ew%�g��g9�e^�yL�aL��^��&���Y�-.kV���
���
�g�,j=]�!�Si>]����k�wx`﬏��(2Ʊ��$J�&0�[������l���o-�p�%3A*v�S���­."��8���g�Zp�U�����f@c@Uq�Lz����Iǎ$6vLw�\dB���zޖ��O�]74`��l���&��$��1pK��(%��H
ȓ�O=K�H��0�	����h+Q��k�woGM�}1^_�;�#�1�T{�^U0�L|���F�ͱ5��V�W�����4P.�";>\L�[���X� >F�ug2��Ͽ�+�	1�B�������𨤀X��tM���_�0h#�J�Z�bN^h��������r�X�,"N}�*F�t�?f
��H�fBj�@��Z���e�>|Q��t訜�0��+Ȁ��H=?_D��u�I2ﳔ��n5?�a�*y3ˉQ\�âi=5s����َW���&�~�4��|�r�0��I��=[�I��Gp�Ğ����ze;��kF/�1�!	����	U�^8䷃�Y���U�Q��C�jKͪ侀;�C��u�7���Vu�,V`��n��
�����nڷ�`�K�֘��)hr��λg�{����`V����))�%߀�3x�\i���cu2oi%`LuՎ"g����v��>�D�)wy����������7�5뭤���9��(��w��ם�4�ݽ��*c�[nrJ��t:21ˌ*��2��C�D����sT5�R�����u:��U����p��+a�pt�k�5σ�^�>�����_H�6��xSph�
@���$�����p�^o˘��3�E�����J�OO��