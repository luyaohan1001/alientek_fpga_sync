��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1M܄>@E�V�(�����o�Ϳ���)��}��]�M,�j�y�0�k��?�Z��=��8o�"���K��;@�H9>�s���]�&%J���Dy��;dO��bi��+onqr�=eng��V�,������ic]�oH���KHn���	��`(�GY��=x�Hj��1���T�Q	S��sgω:�T�14*_[e��GI����˫�|�R�z�:�Dp4	82T����x!��H�뢣�lgaNp;�ؒNǈxpڥ<l�cF�;�쵒MΜL��BE�������/EH��Pk�{zcC��]��?41��$������>��zC��WMæ/�L&��7b�+�}���U/�VB��*��^�/��F���:h1g����$����/�� j��)�]g:n�j8ȈU��G�2��N�3���X{�O��?�1�/P��i����g��LWq|9aZ0y�'Sx�B��2Qe>�2م~�W�a{5��,]>��L{�x��:��P8���L��Y�����.��~���
Q~/p��q �-�=��'��
S���]^��f`6�h�*����7<��ή��N���&���.^X�)��Rcq��է������H�büF����3
ذHV�Ӗ ��J���`ū�������ض� ��t���<�2��d�f^#�����NNi�Ͽ�¹��>O|��
iC�o�YQ^1���CT���Sќn������b��s�~JqƆ>���x��ȸ��@d)�-x�Ӆ&�4���ז�vЪ-�:�����7�� 7�KϢk����j'��Z���غ'���O,��mx[6���]��#���T�9�j(0(#��+\���I��=E3�f��Ⱥl�M���	��8��v�$(������n_֡X�ZqΔ���T�_�Z����D�E�~g���L��ّ���К>���V@�2YW����aPp�}i���� L̉��b~�Zu͕�En��y�1^�����6�\���r����<����� CVD����	� [�g�ǜAL 4[��m�0���3�&:�z�]-�أ�I��pU�i���Ǣ�:�a��#�g�*���o�0��8��Q���	#�6�\=S��O6B9ƿ�:N�-d�
"v: ����&��_]Q.GP�[0ə9P'�OH������[��X�)�-Zv��Ʃ����qjp�U"��Ҡ1�W�qg�`/	x� �[9:�n6[X�nPb�)����"��;X��>~��27פ���Ɨ ysp���R��M�P��O9v���s�93�A<
��k!XD�IQ4�L%��%�MD������f45.��p���C�R�A��(&,�M'4��u�Z(�^k��Й�kk]��>ͬX޽�[dnW{�qT9�-s��l�
$C���1цzW�?�Z�*�u�M��R��k�:��_�j��8�<���O��&©=�����OLtw����َx��_�w��Xȶ1a	1�LT��Ƹ���ޮ�m����Q"�@���3oC�;G�ϗh<q0D	��8�|�i<��dD�Tj��
e����AML5�4�x<^;B��U�o��m����Y;Q����#�������Q�4_b�����d��0�5�&q)Q�֋[�]�J��6�b��G�Eʙ�ܐuy&����H{���
���������\��^�Qٓ�� ���i1�GvC�;�F��MR�q�^RZ}��7O�s��B�f#�j��%�����vC�� ��a�:l��<�m��l��G�D[&V�G��N�`,�@���`��tg��_�^I���{k��<ls���ES�BӐMѸ{\���UL���,�TK�1�_�鮨�~yġ�I�Z�VZ"*ɓBf�2�ب��×�渊F�۱�<�!�22G9�U��@�v��M�R�C�;��2
�w�ue��]*~1�r�W��ש���=����q�T�n��R��b�����;y�t/t��lMt��)�3/ul���,����Lk��s׷1/�K�͈�Ū��ťݿ��y�c)�UfM&�uMY?�w#��́�%T����󕙵��:��c/�����e���S�~�f�_�����jg f��F ��0�#L��9:쓜+�����^�[�t*ҵM�B��y C�g����3�'��Vۇ~o�\�6ʪ�1��Se,/���G}�2F}��X�I���iWҲ�6�o�v�=���ѽK�Z�m��Y�� ���2X�0������ +-�f�:uEɅ��q�U�e��jW�k�sE�5
v�G�a�n>��x�)�
s���C'�8Oz� H��҉8QVA��v��/h"w�����(
��'@���B�6�j	�9i�P!�G�˽�\���L&�����i��Xr�^m�峚���
$����Yj=������e�݈�D|Z������h�8$��c7��8�*�b�ԴY7rCw�B�Y��-����$�]G��j�k'e�ϗ������Xם�f��b�X3X��멼ou�P��(���Kw����_Af�PZ42��uVΚ"{�Hebw���1� `�4V��P�k@]�*�khqL�=��4 Gsg��x�sd��ᄉ �Fm�B�c��-�X���{�vh��{&ޗ�ձ9M����S�F��N�襌 <]���M�F�-1)���v�<���i��g���rp�z��x��t�� ��Z�,C�!�C�7�:j��{�[Z�!������,#��\����ԑ�	��`o���c��m������4t}�`��B|�pI����j�*�k�nM����/��Y��)�>	��.�5\v�[��I��JU�����<��<�p��e�o�u�Y�U��̯KCS��I���|�3C>/hڗ$���Wo�n%�cLd$���v��8<�'��X����-u+�&ޛZ����Zom��c�~����\��O����s9'w`����xo|���*��<q&�5W( Q
�U'i��Kf6v��k�,DQ��q�~	/)DV���N�3��؏�_#�.8�c��0�:��j��;�l/4-`�F�'�X��'�J��
�k��?�{}��~�ӆ�u�+��|���@����Ms"�.m�GF\+�Zx��(�� �rJBM������̇%7j[��s���|�X�K��h��x���:�U6��M����qH�ҡ�����t��-���j/��.$�4$�Bg��,�ω+�o�
��cm�yB�l�c�E
cu�]�^�����w�S9�!�cw�1"&+��9�5�o!?���^pJ�bHP�D�]�������C��yZ=x��(�yr�c���Q���҄�ޙ�Wc�x��2�Z��тm����l!���4�R�:	��iۅ*�ĩ+�+U2~W�eb�U� Q�S��N�w:��=:�)�2�#�h8܃�FpӀ�;��r3�����Q�N�G.n�@�M����.�8;����������I���ր���DV���Ĵ�z�F��Ɍz��.3��LhQ\��>�ӆ�����z�ר��>�Mp���|��3�ڲ�A@3ce���-:��U��&�9�F�K�����O�=��_l ����3�)���nt�*_�'�\B�ck�5X�侻ʃ��+;,u��ԍc�a�Wl\�7��w��ސ���x����^ZY��f�*��nϣ�w����e�RɯA!8$�St/� ���7w���ɥ��܃�X�1U5�ے=ƦQ����!�n�����0���h�J l@h�	9��3�<(�Dp��3���mZ� �R#�T�����)1�)�N]_J�2���_�>HvĶ�,�*mh�4�MF{ K������ǧ�x���
 �{~����Cmi�A�j8.^�A�0��$���2�� �Í��x��<=زy�vR-$$8��e��rҐVW�� -��<�����麹�i��M
4.�?}�랐_���)ymMµ�a����4��dazRw-�)������T�C)�D�݂GX���&!*y@�]�O��9��U�pz��l��{Ob����E�(�6����G-Ubz��� �0@���G���	e������z?q#��9[�F|�B�8*��$/0�[��J���Y��8h�Vs�����F1�%ή&{�~O�[�	�b��Y��T>�W��x���k���bI�w�-��i�>dh��9�k�����4\a��ކ Ry�5߼mF�}s�DQ�8�~�����I~tb+�,��T����,�	�jj�lc)�)6����[�x�bw�/Ǌ�J�ɂ��\�������C�`9�u�.g~|�/�2@v��@0�I%_ 0j�=ل���kTL����2�1��a�iN��x�X��#�
=l�2�ɢ�Acy�](���3�I����,��>��ϙ`70�^5����?�@�ق��:���b5)v<"�����{�f��f6�p=.�C��Dh�@�!>x?�!bQKM��=$�<�6~����>�j0�S���#��|�W�9�8�B����t\��}%�'nv���pIc�
�lŏZѿD�@�0Q=�=���O��ЗP��bf�l5�l���*�.+�N��o������[�	�Ɨ��<)�q�/�EW)��mF[a�D���5N#��1�����@N[����Bv��i	�����	\9@nƷH��"�͖��g���~��l �lY_��m�G��� X�P���S-1�؂0\ưV�4
���r|��D,��Xѭ��p�A��#����|Bp�r�����1.>�q������1�\'Ԓ�w:}ǡ͹��UIQ�PO��������e��z®�QeA�iYؒ�h�C�B���<��s�����>V?I�_M��|'(I�t��	nNP>5���������p����F�]�lJ�L�����i���)�/J���w�v'��}� ����ڔ�9"��:����d��h^L��=�&iE�,��Ļ1Eʣ�ΪqԷ7��=|z�ϵZ��m˭�2�a�Ԯ�Y&��&W��E�:g��������j	��sw-��3���~S}�g��44ß����
���]�[Z�g��J�C��F{!H,���d��WԢ(],��^�E���R�v)�o��R
��U�Ն�C)�����@�N�WQ�Vo���b�1������ i��|=�r�w��G��.F�B��k<���H�O�ul/� ��*��>+$�$���f�j�u��d�iGw��ak?�5�\�ԉv��E=x��-TN]Zt��yչdu;����{�Z����ow�D6V��u��[wW!)|���g�X����F2�r�qx�Cͣ1B����]S�ˤ�mL��g#�|d����0W�B4s��p���N,q+�¹��_j�Y���9NQf�=(K�X
����ް��Biॼ�Otevw�L�Ȣ��PoF:�a���չPP5�k�P~N�C7=�^�/sםW7�`':+����e�����B��l�D�I_�,���X����.#5�zy�A�!U��F�{9��:H ܾ������̬u����&�	��&/�6+����ܳ�8�#���-C\�m}���A7 M�V�g	rw,����*=�:N�)��|"�5�Q�i�:/�>E4Sy�vS��(���xҸU��7�WO�s��U�*�a:]�>��j�<�=�z�-ќ�?�^���09t��������n�{"�����"}�6x���� �'�S	]��C+�X�%�7�:�K�D�c��R�D,�U��xp��h��HWȏ�u=���˓���#Ao��ڏD�- ��t�\�C��Ņ�B�<�J����ڜE-�܏O��Kp����9���C@��z�97���I17h	�jşI5l�`���w��n�t��(ĠBx\"�5M\����d��@")�:EH/��&a�����P����gL�/�˩�*��r�������2��=�M���� �b*d=}����x�~���I�C����2Ϯ]����W8�ד�m�A \\h�a@L��$WI�$<<�@���F�f�gf>���ۼ=�؉����?���Id�Z�����m�W"�{��,����\��W�:Z�	j��"y�2��+2�U��	=�yɿ��҃��Q�e��_Ԃ;H5����d3��3�RH)�(
$���y]�9i���1N˴��eb�7�9BLl%��6�q�O�UǯSC|����KPB���5����I���9�V���w�f��.�)�=����A��\6]|�0�G�9�i$N=�>SD� @�z�Oö�%	��sb ���5�8�t���k�Jxm}�ANr�۽���DV���W+������W���i��4��޺=S�?� a��<7v�U���Y���[z�Ŗ���^.��]`#��I�~���̈��O��VXw�1���1C�}�e멁+}3��Wb�H[`9�v9n���S\�"��p��Ko�F�,	�?�K���cx!���q:bl
"�����R
5L�&@P����̟�P��*.f�h�6�����1n�U�>㿇��,"��f�ȩI��,����c#�|"Zn2���Ii����E��n�6W�46B��kՏ+�]�h@�<�_*ې�<F�c��-��/�R�s�3?���Kdh��ÞFA��u]��dD�B�sX��Mal��y��Ǟ�ׁ�ʔr�	�/%�0��9DJ��H(���h��|Dy�8��z �Պ��u�+�w�˳>�l�AJ++㢛�_������ȣк�k��`W,@>ӣ�"��a���;e �����E#�����MVN̠���g�|�w ���N�=�T��>�z.ܝB���R���jG�����X���IZ��M+�<�2�z0r�L{��rxΈ=<-�
�%0N�W�]�y#R	d��M;8
�	Pi�f��{�(Ҕ c�|~yJ-61�/��f��{)���Z��7~i`=_5�MƱ��Ү3.�WS`̫X�}\/e9�qX�F�\���6�vAD�S�D�J\���`B������T�/D�`�TԤ��0��<*,\3�lI��LF2q5�(p�!�������g<y��~����x��i�Ds�?|�3��i�U	�do�T�CQ,]��{�������q��I��7u!��a��Y��Ss�{�]��o��h�B���˞{���^����TJ��Lxd!�{�|~Rw+��
���R��!��m�~����+��?~(�8��f;c��-sM��[� 4����"�8����by�l�A
cHb)�������A�3v�,/FA�SW���މk��\+]9N�9OX�E�����%B�(����[��]J�[ez	�԰|��5s(� !�E����5<���X�F�i��$��ږ
F�'���]��~0t�˒J�iٔ���S���i
a�`���S����|?����R�yD�����D�%�Ξ�uM؝���Jv���1N��\;*��ƅ�L��(G�p�D'!y��b�X�t�N�!Z�2�S� �D��Z)�t��q��Ә5�%�ߋu���o�g~���ѯ��2v��ڔ��C�~��R��h���~a�je:�7��x��߶-�ԁ�.\�5�B8�F���5�2p��ȥ��G���)J,*q�l�D\ �MCn�XS� �v�'��O�u{PH���= �G���-���`i$:\�����;u9��ZCVd��+٫c�$��$q]��ep��5�l <�q�mz��r��m`i� ���@\�o�\�?#J��*��d����p��]�2oP��ˀ8|��'���>����	�t����b�(�k)���y�L1����������玘�Xb�0�u1���Ԗ�y��q��n��)��B^O���	���)�1P��ot��z~������s�
����n��V���C���������ج1P2܌�4+_��%��Ml����L�h��,� S	A�;�Ӽ8���:�%�VQ�����-��sO�|��\/�\�$v=c�]�AE�D��O�{�l�X���5�%QZ�6/o9{��7z��|�!@�1����a�S� q��ǫ/��L?>>�3T ���1�"�c�w�T-+C�;��-��������ȶ�z^���C�\$�p>���(���:��������|s²EO(�3��J��b4hN�QQ?�ҳ�.4p��ׇ<���V�0|ġ�SP���d���IP�����<۲��r�ب��y��8�+.�H�zf�M��`���a��P�O�*�1Tk����u^��=�C޽I�౫�?������_��3�YcF����mM�5�u�>s3@$�w����5;ҍQd�<�)�j��Xs���\u�����6�٠��z���F��9c�M%���p[�s4�mU��B_g�d���%�������!�u�ZΨD��Y�
�;7�OL�y���B�M���,M�K�oz�i:
��;�;�aM �w��|���IBB��t!�L)�c��,�M�=p'I�H�"'?A����gJ!&���-�bG��&d���l�`"������� $�c'�@�K��� ���'M	����k���<�$��<*N�/P�'��㧘�ó���_�'�Ԟ�(����r�*�&jX�V�Ű��j�Wϓ��i��w�i�����:�M�1�h<Ƙ���&�l̞�(�����h���LA�+i|71I��7��<Lg�	+�,���X�p��4!��z��P�λ��]wDB}w��ȥĶ�=I,SUP`v0��I�q>p�8X9?z���&�u^�6�����ێr�.��*V�2�a�&�����3*H�:3s �I�� q��Q����	@Ի+LH�8Wz�c�q��e>��ϐ�&���u@�輕� iޞ�J�dݸ�m\�ބfh�kY8s��� Z�]S���~n�}�H���RDP耮�l��s2�uŸ��kRF'NU���k���*m�i�{꤀�����N�ȣ'ڽ�������*�Ƹ�Z!ـ�߭��.d���Xq�Ta�XO���A��S��
e��K��Ze�Z����5h��k,Adu�\U@�����`Y��p�*�KcW<s�<P<����.C�Z���#:*;�~Is�ꂙii���J������ 9�T���	h��<Ĕ2Bc��2�n�ɽ�{e�JL� {:݇���
����1>�Fvf׎2`������	�	 ј�sۆ����]���.N��s$9;g�0ar�� d�w��Ol'����`[ZQ*�2����(�0�6�@�+��߄��9�: 1��e��܋i*�0�1���g�m["��5$18�K:h��S�X<��K$T�ϸM�8��n�Y�3x��܏S��W�e���zʧ7�n�Yk@곉��T��ч�t}�wQ�y̢m�ѓL����x Mh	��M�	h4fn!5��ǌ!+�-��ɫ�o$�&,�!%�@=���� ��=7>�wo��Ղ⇽��>�{0�J�n�/����4�����^W��L-Df^�0��LT'GNb�t�I1H3�%��(��"$`#������a%eF��P;漏 8r��E}�cL(E��}_)��]Hr���P$��P�AR�>[,� ��ժA6_"?��s�l���K�{ ���׺"��->�������e�g��{�T�,�v�]u|_TН�P/���g����"����5�0Z ���ˠ�?�$C�
�/��)rZ��ղ�f��xpތ��F�?̹Փw98[���a�����bfW׹�2�`�E΅��*sZY��d��-(9uD4)�k	��0!�-vIQI��C<�������A�W�h�-&Q�d����2&x��Kt��Mחơ�-�Ľ���{����Z? nj�,���
�	�_������S�;��cH���+���ԫ�4��� ����Y��CV<P�ga~5x��A�Ao6R�,�|���|q[4�o]�����V�g��KO�g#@�Q���6�]���V��oAE3_,۽��/.��%F�Lӊ�"s�=���R]�x�"�0~��Y	L�30��п#��m��]JR��q�0���+�h*|3� ���駶���xe������������!��	b�>:3��EP+xH���>7�[%��d�g�Ѝ�i���u7�/��f����b8�H�K�/�G�祂��S:��R1��qmTLza��A.�0�c׃���|��w�ۺ���2D'CW��ۣ1�U�6[[�pM"�g�_��'4�_ίC⛧>�����cc��f�w�����I�样C���H�N� �f�#�+Շ׷9�~a(k&�~��.Y ��{Ny�Y�Zy��;$����N��t�F��#�qm�J����ڬo��sX�|�jq���K*�n��Al$�����;N؂<���%��V��s�}S�u�e����C��b�I)�4.��;9Q�凮��iC̀G�%�|�Q�W��1�5��H�$_�ss!:)Cw�[�SMX��JG��D�6h�&-�R����pMH�c)T�>�����I86���N�Č��#͉mO<}�i�J^	;��U��uS0vJ���;ç��|Y�j`6��ۆ"�H���}������h{��vX�i��&:漮c��]Ҽ�Y"��x��o�è��������,L�iñ<�/LG`r��b�����WǷ�Õ���kl
\X[�O����d�﮷��/��je�Һù���%%��L���&�>#�3��8�q����'�8�����q�2��h;�<^�^����.ѓ�w\s���v8�$::�}?;���H�� �����<�2� qQ���Ãè�y��؈읠q� ���H��G����2�:R}P.D ���6t�c���ykfb��� �.m��`3��bO>T1�E��-$]qL��j�ZJ��h�T�����]��7|�����t^U�����g��(EG�� ���[�d"G��aYOR������7�(����>.=��z���i֜�y���3����4���/F�VPA��"���=��і��;t�D��{��4(܊�^5�GydQK���?��&�8�����ʀAA�O�`m��<�(��C��<S�TaNZ�m�Y�dO-h�ͷ?P������b<����mYoۋf3_���2�x���tj�3��6*�坟�U�sm7Zj�=����v��\&�,�߬-^�B� g�Zf,R&��$��M��[��O�)ĕxzCO��//G�{�'(������	�ѯe��4�5���wJwr�T+M������5�&e��j[	Æ��b�9;�3�R���D��DQ���*B�$;����ʖ��U�c��<�P��ѱ��@#�ôD����`{�B���l뱀���&r�}܂�B���	vb�B'�	)���	&T���:�d~G�Y�*��C&��]�m~3�����V���m_�0�17�6jl|v�m�!����G#+Z'������y�#�m_�a/]��iA�1�� NZ=W[�sN@�{����dW#F@ߕot�#Cv�����T*L�i�4�B1��j��]"�5Y��B��b����V�e���a��v�h,%^M�l�"�`z�,YK�)Zt��E8����B�e��@�����l�M9s
�j�����o���~θ9S�k�xE0��<OD淈��s�;6D�u�U�NS"k�[,=o.�����ɵ�H��V���
-yq:ǈ��P�B�K��敥�`U��4��6N������h��0ub|�JI,)F@�y(��c~=K�9x�DmM�S�(��AS
R[d"�e�z�m�&;I����%�rW�-B���uP�����x1Oq���S�H��ٖ����+cQ�Kځ(�V~��������{	-~8�2E�H�(��)�g�/��`_��wH�l�	�͑o�bn���
�^��!��ׇ�tl�=Nn���;�!ܗ�؂���}��u��(��6f��V+
h���ZoTq��6Ώ���!u�V,�g�Bh��pȗEf'�� ���D�U��?�Z84u%de�O�I�D�u�=M�5*��J����W*��d�8�͝x;�g<Rv�� �6�*��LѥD�Ƣ<��O�Њ� ���k����q�b4���_(����Z��-O;t��R��������Υ�B}�]�p�vW�o&EyG�(B���,���j>Χ��۹�T�Dn?�-��+;��~��k��=���ў�e=X�Y�����L��d����r�e#k�'Es#�5����@pَl�	�+�ᤌlP�@ް���2lp����.�q3��1j�p���F���k0/c2i����`��B�Q�ea�Ŗ���lR/���b{h����wPw?0���3ό��x �o����`i�K��ۊn\�8e8�p�d9{T��	�=��+��ɗ���s0����<|�ݦP,r�բ!0�>�;2�u(=�>�b���?�E� d�<�p�V0�Ÿ����18�6Ib�����v�\o̾���T�:����᰸F����Z*	��I)|��ǳy[�La�H{8΃��.�׍�?f���u���׌���@[e���d�c񯢍�� ��w�K���r~�^���J.M��,&��)7~t���$��{c/�p����~��y�W��*��9!i��d��͡�T�ľݪ��OA�CF	�2/��U�ш9F#D�sޓ�]3"K9p��,�eY}�15���xj�⏉e?e�;U������Mow���z�[a���\3���ET���L�.YC�ơn�(My����3�=8;��c�N�ji东EBV=��7S,��q��/��QvU^#4i�=^8f��xx��"4h ��|J�׵[q�H�~.�j�a&pz�۪'����ݙ�d�	c�q����RJ�������>5O%������#c/���崓D�Nັ��7��/�ka��L���"*���t�/�oB?�'4�p?��|���Ltd�?z�s��{����ée�f ��K>a�	t	�W������HH*D�}%�Mn��򪂌��a%¿�{E�W�N{Z��(-Ar�!�q�~��(��]��7Ya�����E׏�f|�-d$��� �N2���������}/N�* ����*dX+-�z�J��*r��g�-�=\�Ågv�ZU��?���\n�k_�֭~Iϊ!Bw0����֧��ڤ~���������n���i�.,�yog/E�٬E�f�.q|JxB!~t5_��F��Y�Ѿ<!���]_�!r���3_�`���0W�	�O��K���|�����×D}����x�A�>BPfҊo*��_�s����E��׉��'�Xt�����L,�?A�آ�+�Z"J!�1{"���SW�O�������G����
���fgj#Ƕ�m���92�1�S��Q�f�34hEu"�s�M|�X�ZTuA+��G���j
��av�Ag�9׳L2��R�x���`��A��r�5��q�k�94��&j��1�$���Z�� <��ԕ@���9c$�r̋\jS$V�C�����Y0�J�<V('�m�x��`l��\��~Ys�IZ�'v��F��� �2{/f�Y�3h��?tE�z@�e]�αN���BF�۔۞W��Y`{�-��Se8�^���4>P��W�Wb~i!j:�C0�y6F���D�IG�Z���s�i���R��0S��A=i�س��R�G�jU^A�(Ƞ�J?s����rN�g�a�n��ʅ�$���WZ�T�p��F9ʓ	��$��hFz�N�j��W3TK��n�^�x��b��kS���W).i�������0��k=}N�,��07ǫm;0qc�vR�+_�ی�=�OS��^5� z)�E�wO� ���h;�g���	Ë\
>-Β;"�:y�D��zߟ,�����Ջ���2"����3�7O���t+X`�᥺�$ܶΊ��W\.�D�ީ����������B��l�o��93�Q�>�n��\�L�	��SJ�Ϻ��^�v�b�Mxʋ��sW��#����=�����̀��RxK*~��u�
��#!R�\B��?�sZx����J|�g��ӓ�	Fq�Oi�&���S�g%�^h���Xk������Z�,`�t9 ��σ+��̳��C�N�y��u"�r���Z�p:�X+��!���=~�$\^F��٘�?Θ���I\����ؕぞdIp�"3�|gCq���W�t�<�j�#ċ�4��.>5��1Č�,ہ֪:�m�U�����-�������R�>T�tە$���������CW��D�f�I�az_���s��4�G���-iXA.�ӽ�ޥf);>+f��W=ԧ�����M�`l�V/=4g@dmY�����Q��T��� z}�g��+/��ucؿ�3�Z[H�%�vM]�<E~��Ol�S�Gx,M��\$3�W���'9+����������n�*��مhd=F�j�L�r���y58�g�f��0�z�#�ߤ�{����2�G�~K����E�*y��� ��%�A+e�"�6]2K�j�S�Z͓x��bB��K���mt_�o�*<#@�6�3E��&<pGo#��ob���� �wF��fj��P�67;����u-'�9ȟ�
���ZQoX߸�i�)VP���+ĉ�������g��V��w��z����Y��w4Xn�o�������~�B�\kP&�k4yR�ˢj%�r!g"{!����x�j��W���嫂�|!���s���s?h�޵�(b���uYN\ŅH.�:���˶�rB��V�bxʂ�'�2K30x�"x�n�4+�ej�a+����w ��[N��V�=X�	[A��n���)���;�Д�A��s�'0�P��˝>8'�����wH�i�j�Upp_>�u��T�th~�#�A6�֭x��o݇��7 '�����ZB��Y�%�#������s2�  �l���7���dS���vh����+��Bqd@����Al�=�������g�ĺ�Q����Y�[NkB��&�&{��K�'"M�%��D5�m��.zZ|��5��VND^�(�z�%(���)�^
�G�3� ;��>TQh�b�$��x��9H3�0�#n�;����Ԓ�μ��b��A Clp�}�'˷��;Z�gW�	%�
���]_�	T +A�`t��%Wz�τ-'���
7c��bY�ǲ��y=��lO��g��;Hg�t)��G3�� ���$Q�-;I<*g+�zW�@����>"c��8����l�>��os�qZIp��b�C�� Y5	ϣԆ��@+����	C O�)�����%}7�V�m�XF�0��9�"#sIB��d��{=�"�vF�>�&��}��1���A9c�ķ�(R��7~��a#��)I�����:{�6M{6p��ܻ�瘝�G�:L���t��J�*[��@oi���	�\?v���5&�FWz��P�m�����LǇ�������ӤfI2i�YgY㔧mf�IC����K�q9�\���Q�����an���HG������{�o�2�I� xL�e��g��9y�2-�P`6�h�l���Zz]�]�*l!/Fh����jr0�ީ��$wU��wj�HW��%�S�Kpk�F��S-��� uB㴸�{���<wԃ�c{Gq:�J��r3��a&;���XeR�ܭ��}����i��e���蕎���(�T������ώ�&Ab?��]X��ŷ8sW���V#��l�Iy�Y��RV�����%)1�
&Q��׀ȏ��F�X@���Ms�Ժ2�ix5�z{E$��j�]jȎ�������A��H����"�W/6�&a�2k�A��]��������#y_ͺ���B��^"����8���&�[g뜵O�x3#ol��!�0�"A�<�h.�{ɸ��S�P��ߊ�@OC��Fϰr&q�E1(K<n�t���S��1սZ�'Bt�9�2��A�隸Q�0��3גK&��o=�KTk�E<��3x�5���B-����q���r]��*:R��$����C���4��+ '���`K��,��� P�pΣƃ�wp��j����ͷ�er�,�o����t�fʸH�����R�-c�����0�����aQ«F#$���j7��79��]:j<���.��z�������J=nd�]�m��;�w���`�K�d!��[l������u�i1T3�D�}"P#t����b� $���q��}�9�+�8lT�|ѯy�ˬ�k2zp)]��m����I:@�E���<��3����{5z�i��� 5��s��F���� �/�u�5�(�6����#��XΫ��8f$ް�b���)s �u�w)��To-P��i����
B�����1�����57أz����S.}^,���#���0Kv�2��o���w�7�3�Q����7A֣}}&��o�i���&5wcb����m�MTsՒ �+�=���:T*�vx��3m�4��Q�U�' � gs�xY�S"�;�MqIzw��J�XX��2��;�A�?���>�Wd4��>,��}_�.��eF��eW�XT�7x��,2�,tiYϧ9����K�kʌ}K�hz�<f���{����-g�����# 8�Y���[��^������̌>���E�~q����s���3��wj��V�9;p��}l�4�XRε�1�4��������q)��v�67�*�,����D���0�z��͜�R�D!�oG��*	�O4z��l�M@uwO lߠ���a�X��Y�i��39���~^_E_ۭȻeJ����:.F�nr���Xk�*;�$EN�6]�����g<!�J#i]�T�z7�Z��#c�E=o��7^=ؔ���B&�N�iGZ���y�9ۜ���aq�f�4�]��j9{�Y����kn\�2�uB�pP�ĳo�Ms���^7�*��1��I��ՈTf}���[$�h��?`4B�9����n�K��y@F�z|G%�����]*r=�,��V�K�[ܞ����2�cBֿ�r(i^��1��{�2R���A�^ sgG �K�݇aQ���B���Vn*I�F�Z�.^������riU��&z���oY�G��R���NI�ȋ_�/)i�ɐ�!	Q/)�	�&�~)3j�x����߹��Q향��a���C����2Z��:��x���@*�j2n����Z�To��dv�,2�손-����)h2#'Ǧ[���Y�Է����2�#�A5-�������3����<�Ĺ3h������F����+����䉿K�	[n�9X�r� H=[չ��U��ZC�G����װ械p0&�(�! �E>����B�4L��}����B��pb�k��[s�E�dX0#{�QF���b�*n���F�,m���P_[H�����.����R�ı�@�Z�ʗj�ALG��ce�,��	|�y���=�ë��<���~��S�t�=�>�҉y�3�ᒀ� t��Y�\s�>v����\�r�t��#�h����,#b��Ohux6�~j�;��{+��GHl���9���ϱ�1��EݬqV^n����01�z?��f��*���Z�������
��k=���ԩ/nj���}�6������.	;���|*U����Nd?Ҳ1Q�U۪������cOhߖ��SlKL���R�1�e\��XW%�`&:�j�Ež�o�+�u��z䎩�����p��ͧ%MH>�q9���6���`d�D݇�H]Pe�l��(f��5��ډsIK ՟����@��]!V���%!m
� �n�d�{��	��9����ҭ���=�J����
ehd�6F�p�T��N*��%�c呻ijG�lg�ii~ǿF&'�@�,��2����"�h�
4d�@��&�.�Wc��f�Ұ�摅L���|-M���q�J~�J��a�A��*ul߄X������f4�oz���?�gdV �R� �&߫��Z��`�nx�����Dc]�_'���_2��
�<:䗽�0���V>|w�������F�;��6����F�)�N:�W��K�5��0N��9H4�n_@�)�$��N��x�w$�~� U޲������UD/�����@���U�6e*>����,��� ��cO����Mb�z� ����	�~+���3'p�ˏ`�f ��}�<L{���7o���n���\bܮ���h��Hx����A�!��L�a6�/��v&^z�߄p��#(��]�[��8GJ�5qj��@�z���n�XG�3�_���
��ţ�o��{�#�b��XW�P���%7���W�%Qx�Y�V(*�����t�@��7���Y2n�sW5��9ů #�v���@��A�jM����*Hf{<<e(\[FFr��8乊G �}�Ȼ# ���EK9ľ�HN�U�'����ܘ\Q��P�Zu0��F���S@Y42����/��p�]S+��M��iXA�:gZ'J+Ι6d)= �>�j��=�=<��	�]�\ !Rv>p��D�������� �(�!`~.�=
�B0|V��7�ζ�M�������2:&�'H.�ng�hr�jK���|A����q�~__x#��3�z� bAE��c
n:.H�x����}��4>J��a����#�`��&�֘�<�'ۇE�?�<�6~�X}��{D6>���d��}�Z�0?�v�'aE@�Ǡ�P�9����=�`�����Q��1w�`rO�QFܗ�.ɴql!�;�#�����̼H�w3� ���^��N��&����G��z��
|7ow�Q?D��w^Nׅ �%����zN4�xF�j�o�ɥ�BL������X�&AdyO)�d[Ցn�<((M���:���^A����o���;P=�^Ԩ���Am%]z�u���N���5��]���F�;��rO�y���)�������K�����z�@���K瘽YAꠢ�����,��L���#�����ض���X.��-1���U
��i��x�qʾ�84�l([l���޳���������s��P���"��Ĝ.�0ظ�`'שy[�VϡS^�a��\ѲRf�ߢri�g�y��0޸���&F/��1Z�j�y�̩'�.�c���$��� ��ܙ���B������I�l�O	ؿ�m��j9���ܫ�ꙃ4C�ɣ�� u����n�)��B����q�Ua�)PY˾�45x��9)�#�*M��	��a��~����K��>�$��D���pǦ��Q������J�,x��M�<��S�h��D�k��#��k�=��V���<�Y�B�A�u�L�|�w�*Q��N�d� D�C[������s�
�Āa8�6^G�%U0��;#�˗�����b��Ѩg薨�B���!�#n����Ȣ!���}��h���\�$xI[�fFJ�:�sx�鸪���~Hf��ωQ�	Ǩ�^S�`t��FM*�召B����*V�s"\�~N��=�5ǀ�d�y��"�nT�Q�J�;	�	hSFP��c�v%�1�H ��d�@v�ӌ4�0���/�{2	#)t1K@s��d��t���v!�Q��}'�VK;�����[�Lz��;{L�2��H����'O�cg�\+��YL�O��P&*LS
���]��Jj߷h��~Ƅ�[j6E} ws��Ӈn�����۲�e�D G�N�qi�ltѫn��S�=g��hd���zJ"�g]�T�������w:I :�8��؋o&k�l(���P?�B����vk���.=�؄�A����3X��{L[u�r���y��)o��&�����z#�e�����I�MK8Әy���'�sC�� C����TyĹ��B&Q������;�FW�~gk��S�PiF��zGI�]��cb������͕��T�>7K䰞ݘ�� �J�&��%�=`:�ߵ_�Z�6����M淳+� �E��\8���RAJ���d�����b������Q%�`�m��Y���`P�sX.r��Q���X�A�M"�.��A�wj�д�-����ǕԘ��ȾEv�\�Xs�VoR>N#���+H��ĦYwK�lvg�H���L,Kع��j~��e^�l����V�vI��Ï����a��sI>��%��*��EEc�JW_Jҗ*!jQ2�����D��z8 ��*��:������c��e}���{��Y8Y��܃���"?�>����ސ�4�����	�`�W4�����9_ΎX{�D�k��	�}@h;%O3	3"��3~�/�������Ms*���-%[�����L���@�SO��A�m��\�����������&���^J�ӂ�t�H���QH���X6y:b)G�݊�Nn�c��IϼI��E�� �?��a����6_+��;=3��� n�C�Z�B�EΕ"v��r�!	��9��m�;�3IV�.�n�Zz�����2��H�[�h�451�M"Sh�p(�����樳.���ж�y����(��ǰ�٨j��~ч\=T#Yݽ�֛,(�|-'ֽyfw^|/�ˁ݅�%���{�J��d�)��Y)t�U�*j��n���D�ˍ�䜍]�͠oǴ�$���5��\��r�q'=��ZM�Tt�������\��x��g��F����ö�$B1����� ��1��}���4v2��L�	G�X%�O�	۫Y�E��Ԕ)��-1?����AW�]�P�I+H�8|�Ъ� S	*�:s��Z�����i�Ѵ]�w6�cRO
���\���(u.��(Ҝ'ߵH��MTQM�H�C�N����* �ҥ���Z���4�]���������������������C�b[��)j;�%B��Gˬʤ�0�e�}�_�k������l���m�ԹD�Ģ'2��{�]�%��`?^��.RYy��i9me��_�a���*P��ߔ�B,�-�i��e܎�X��(��9c%���kynʭ-5�WD@2Y�+�D�C+&�
{�2��HIy��D2A��&�=u����Gov���L\�鍃bl�����7�E.^I���w���ޫ��K�p��oB"���0�Z6���i�?�E�����l�9t�J�]sJX\�m��nJ@�Z�/��t��m�M]8X���_RC�@��wϝ��8Cv�Q!��</+�m;����v��fwejV=�5Sݽ�s/ѣ�@�*�w���γ*� >{�0Oxw�>�����r�{�dU`�P�m�xrT�c��je`p(�g�駮�v����t؞�p:b8���!K�,�[ʖ}���hP�6�]OO��&��b����jQ���!��,
Q&Q�_=�My��Q���]$�(/�g^�W<ud2���״�!��v��K�\��r�R��0t8U�;P<&�@���G�7�fpmMO�v�{�.g*ֿm,x<����ڌFU�`e�Iѝ1�`�,��8�S�Y3b��Xt#fy>�c9�w�az~�Ĩ�ܮ�����%�֗�n�o��CS�PmW& ��˂Ū�/�Ik(-�aN�4͒������& ,2��t� P/y�㪤},��
d�hj#2g��T
�l�{�^��
��3
e��M7NC�^����L���
�?mF��ޛ��tY�@�>g���6H���Ѷ9Xp%�L�*e��{����o��ÿ�5�B���fg�sD�����Q�G {���_�G�%�r��Pzo���t��'�;|��7>���%���&^�ؾ��?�[��`�����ͳ������G���-��Ç�{��E�7Q��l�&�$m։F�`^}YHj^����.p2��F%y4���n'k%�1��D0K���t��3���(?1�Y��`����&�:��W�(���RT<jz"y|S :�bh�Yu��;�H8ce��1x�s�q��ڍ��u���K�G[����؁[��+��=�}�Fj��������8�=Zd��a��y�&  "ݕ�j���4��#��bt����;N5P��}��w��t��8�+��e����t�ĺ���@A�G֛.�3�+�	����CK�[�yiߨ��s?-���A�������7�RܼD��(Ե�\��/�1v��s�d���o���a*<u!��#��֪�����Z�N�����G׆.�&~1�"ƻO_E�*�"��N#�N.� +�,�0�H�#0���%%�ʆ�����=��p��x�Z��{}_��578�[���q�C;�M��I�8�!)&�8�p8�W �3�jH�'����V4�
��L��`8/e	��1�p�S�&�t�r�oD�|1��lZ!�n6�����(�p�����O���Nu��Ҽ�l�Cnյ�a�1q�,Ž�u����(��;����"����⟕�=�wH �*Q�;����C9
ZM�=���mi�V����Zc��3Z��!î��-7����Gͫ�p����P�2t�2�,mi?.I���ޖ���Zk�����!�����ӓ�b��<�i�r��m��=ʞ���σ�0��Un�I������~]�Գ�c�[�ű��:_�o�݅~���d�
$D���:��a���~:5���v'N%�Q�ե�OF��_��A�`nӟ�?�J�xr��J.���"������J��@$L�r���2]"]�Mƃ����7�m���A�<�VV������3�`Ok{]�yg�*�@��f�s����Rh(x�4w�q	T���3�-�����-���,�8���/�MO/��>Z=y��<���u
X�SU}���F�F�-��g�U�(������H�F���r^�.+L�{�$��P W!I1�9�K��cК�pͼ �c��o��G�my�h�?7A���)"����o+����UַpOML#�DEn����ExB�浳�L�[�"�|Z�A�Ӝ���ղ����*����9��E�ХPsX�h �і-���OJ�K�����EljsO�X�c�H�!^<�m(��^s?��b>I���g�;dyi�"6hL�p���}i�E��%�K8G��je�JRjDFإx�%�[���s�j���rՇ�h�M���7-ԝ��k~���k߻�5�H��r�K$�Fۦf�a�T�B��H2�Y�a-�������l]�0q|Fh��y���D�ٟ,<š㜤��2��25~�I%ɔۨp+���9��J�!�Q��`���8���7�W��4t����Y���.�a����8�r�$�齻���F��S�3�n�h��NP���+��KcB��x8��1�NU_L�z����Ί�v�6�����ٔG}2��Si�d��o)����w� ����ΓU�]�^���GR��]�&�P6��?ҭ�LY��$�,�|�I욥�]��֓�s[����4�A���.�Ӂ;���Ժ�]�(72W2��5B� �G��ٽ�f���n��S�!p.e[f�<�ӱ�sp6j�10	�/���|@ѭ���N�x�H(�=�!��,��y�6���|�?)D�X.�m�/OuX��˰�Q�c�m�z2QFnϗ� ���8Ioa�$ϐ���(Ml� �EW���`��l�8PE�q-j�xE�7Gc�O�ف�<�����i��&�������=(o~�9�+���$�H����b�D�"'n�&���Xm)���)�=X6b�~�M?��X��vk��E�Sϼh����-U �5a�!E�	o����}���k�(����q�:6|��m�$��$����x�۽F
�Q�!Z#F�|�KwI�����hV����x�ϓ��V���)�5��ϓֽ�qI㙷�s��p܅�t������~U�Ϋ�ϒq���37K�*z_:)�j���{7"`�0\9���,��3 a��ӗ�A�){'�� �f�c����Mҭ5�wDF�3n��t�n��1��
�L+���]�p�]m�����9M�0��S��}�I����і%!|���&W:쪅��n��qqE����ۋm��PCۏ`Z���E�#� (���P�����T�t$�_O?�5���p�فP�i�k�[�0�⟱e�Ћ1SQ �D��Cv'҅3�B�g�O��wr��u���^�}�{��x�\4��Y��}	Dy1()�VU��>����(y��R���v���e6)�;��{z�HP��<>ט���G1F�볒'�#�P���{��ݜ$�".�H���e4���~�En�������,�!����l%AR���<�>OMߏ��W�+:���?T����79�@Z��vs�sA e��쮃�e4��	Zv���8��r/X����d�,#8	�bU��]'�<�a�q�&�''���G�ِ6'�oa������s���^W- tQ?��@E�y���l��I�OB�p����V�D#i9��[�F�y���O1(��G�b[m7
��ߦ��2k���TB�Uz{�����;��� o�IݝG&$e,S��f*#P��'xq�pfS��r�u�~y�$� �]�O ���ڮ7y٬wm�2���_����-������N(��E�6��e�U�hS��Ar w	guTI#�m_Ҩ7^EB"��H*�4���ϼ<Aj���RqQ6:���b�Pi�͖��_�R��OP�|@���m �$�P�S�i�U�A;�|EVx�;x -�bSU-,jP�2�`J�n`tg���p6�3�gEf�.���rF{:�!g8�<�]�v�Cc:�eZ-U�3{($hg�J�ʔ�D���\�Y���i�KF���~"��~��\��i����1@`b�:��3�'���_��=��������u�x<��w��~��`�6��N�R�qǼ/�M�Y�2U
�ۓ���籦|�;�()p!�k8cE�1���:����I�US0K�n"8�>ޕu�4� �ϒ�o^�b���-Y��><e��fB���}}#p�T�I����� .lg��l�_a��(G��{��o�4#�$e5���5˚#�b�I�	u�m�ތ�	X(�յh_��u����zF�]��x���[tZh�Q�0ZƷo_����Gz6)7|�aEe�~`�x�Yk��<\j�L����N3�t�;=�v\�pͪ�NF�siB�ēq��N����h��G�����g���-=�݂P����,2�g�]��r�2U&�lB컭`كa��v�R��Di��,a\(�2^��]b�iߠ������ot��g��_]5�D��C��`!�[հ�A���Z��@�s�ݦ_�A�w8=,yp����kX�yם"�n�j `t��%�V� G�x9�T��dD���r�\1�~�JP��J9�ܺ���A�Yv�c�(s�?{ޣ�7E��|/���|y��r���9mi%F'�����%�^KH�9��������{���"����6Ǐj+,F���r���0�}�?5�v�&u��'#�����g%�c��tn��.En�2V�k߄��y��V������,��G4���,X���8;�?i1�!,�'��ʺ�<բ$�I3֚����1��Ә_�����Q �2����ʅ��1���v�͈В?	5m���۶5�4��[W�?�5��Z!ܹ���X�t���O�o� ~���'����H��|�^2Ҩ�	�rF5�ܞ�̱~���f2y7&S<A=ĿG�k��{�&M9n(�+�}?|z�aͥbI �XhV�6L;���Hc��|��:����c�'�Z#�pˑd��l'�����ӻq�oy��Y��{����4dDF�F�6�o�!�8�~Mh�,�P��=A�Rvs��B�Eomu�lT��d��3�S�U���n�BA�^pG�����ّ����w��q�q�@�M-�� +��j�{�dj�Yirr����j]�ȍ����-��MT�q��fDvt��-�r����z��W��(���Ѱx����2�@�����_�׬N�MU���ݘ���2�!4 ݚ��� [�H��W�oR�̆VD�H�yX��_1Q�Ju���������Z���IvLХ�.\��A��w�j0#�I
f*(#M�� v7�)��_��[�^w_oH��%SuF&ܢ��?j��Z��ɞ�TYȝ a`�"ߺ����h�͌�X?��m�T��20_�Pt�Q#}^5 ](�px/}�9���C��qq�X~�n[�����Tj�B;�����u��|����g�컀�*p֗�˿uN�Tn]�j�?������t�Xo�P���T�y�c�Y�%G?���=�[8~�۳���&�����!�j���e<}�CtAxB۞�by��Y���T\E�6A^y��O2qxb���.I/�kͥ�H:{/���[.��r�xOA+f8c�Kj����$��C<)�2�b!y 9z(��]�{"����d�������lE��aۓf�Ɲ�\��.�F���l"*�3=�L	��m��t����ڻ�6̿+��5X�ڻ�Q8�ɏ�������@�u�$�k��R�V��[�Ƨ�
�'������yJϞ���-f/���F�ʥGg��͠���N�+2����h���u��c٠��*g�2�_� �%>�9x�oO��/lL#$���2QV��Jd�E/�H霝����N���^	�+�AV�q�P��I�s���58�x�K�Մ��������R?B�e�󽋳*�����%kr�Q��y��~d�R�4L�)����M�$�N�#��G���Θ�J{�ܦP]�����~%1z�T5��u�e�F�M߽�������:��N[&�n��e*�|�-]ZM��?k3Ds�yu�ˌY�p�H�������P��J�BL��4�1��?bC��oQ m�&�s'��6��7Z�p�>��.U�g�&諔s���,X���e>��cf�N&V����#�q8m�m���E�Y�z&�����&%�f��艂hˍ���P�akRq�%f&S;J�Y���@�D��i����'@�
ahٓD��ޘ����ێ�|UM!�㍈����I%�hs���F��6�vC����EsHY��6� �ik�� ���l����B)�8!�I��=�'Jo��T��S�;Zm(�7)�խ��pTv�n!������7$���W��X%'���G�+kR��� ��+��Y�a�l�ru�*`���d�D$R��"�����:�q��+���T�i�����$��9��1��	�̢],W ��9��]���C�����ڎ�^em8�v���A�cD� �Mv
_:Z���}R ��8@�C�덬s�a��P6�$�#�oU�1�?x��w��Q[���x����i�_�}ؖ%�PE��<:ԀZ:N5�0�j�aD>��%+��)�қ%\s��At	��4-�w̡0�ƔvAP1ă�'n؋I��S,D!�4��!4��`��bێ��#Z�3�U]p1ܝ�خ>�߹�U����Sg|.fL>c#�����~���/�}�~�b&
n����qk����?U�K;4:�֮S��㶛`��E,f�@�+�$ByHG����`j!r����ÓCCZ�G ��@�샰����h�'��5j����և�A�%��~1 �%N/�ʦv)c)S~al�x��ܖ��~��O����1.���q"�H͛��9�
��a��!���0%�֋7���O�h�>�N9�Ck�Qhwr�;a2�s�>GJ��=�qz�u��T�%3k-����ۢ�p{���oI2Ѥ/��ޯѴ��.o��?zj�x�?W'�4���J�u��Q�+ꇪ�s��/f�|>���U��1Ԋ�W�˟���g��S�O�����þ�#R��l_&�Ԗ��,��Z5s��A�WO'��S@�dl�O����[S~.�(2����}�I�	WjWm�������{�s����o��t�7i�uǭ���V,�[��^�����ĭq�g)��rJ��t&{��f6������b��%���������U�4��W9g�N����tz-�,%���8��d|���4�_�($�w��@�ҳ@�{���\��k�T�`����DH]�}�Di5����Ǯł�mKTct���<m"ߨ�۲��x�=�挐���c)��\�l�x���F�'!�ٴ3� \U�U�1�%�o����"b0t�<b^e���㍟��s{�� ?�2�R��=�N`��)O� �A�be&�1������yۮZleN�0��\�T�y�Q�Q�o�_9����Cg����p(�������/V ʪ�@��g�"���Zr��G:�9��.�8*������
{xy� K���I�d�d�Ƥ%O��t�g̝>M�l����Ga��Z�ʕ~I32�?eti���Aւ�Χ1t�����y~5~սYV��CfK���.1I�%c3Ԩ6PA�7P<�"�4��>����%�G�S˥����n�����U��������DMa1������nã^� �v!�tG* j� �V�ċ\f�KӴ78�����&�^`!P$�6Y�Z��z����ˉ�g�ۚ贁���KӍ)�U�d9h�F�9�u�(��eU�����
DLz��Q/tX!�m%z�G����u���_İH��r��Sp�AH�9,#�m��V��BzV�U@��Ͼ$o�:<i�@����)*^x���������x��O`9�
ů�Y��%�!�-�(�ᑽ�AA}�K��E��P x��ѝ�� â�jg$���@d�]����Hifm�O7ֻ���#�Tʧ#\��A��6��e�0�g���ձgn������������S$�
ɷd�j6���M�{�>��[X�0B�k]��O$��$�S}�z��l�+y��(�G3�r@����f�A��[�*�$��W�({���޹)Q��=4���ި0�~�R����&����g���+��<�I��ɐ�Q��0Ak�cu}��3��2p|�-���'.��x&�L���Y��4ytU�H�5tC�G�d��^zl;r���k��,L���W!�.����d�|�<�w�+ӧ,k�k���N����Qf=p/�jtd{3����/Z��y�_�.gߞ'��r"��7c��I�H/�I�d�\����RY��Ɇ�x��4Y�r{Q3�`719���4�=�:��M��BǬ���R�*��k*��`�����-Ù�h���f��fU�V�V�T: \��I+L�4}=�IE}�� W"���c���YN'{����Ǻ*���`�� ������4����3(�@�%5�L�?C�R@�ܕ:G+$�<kM�|&3����> r�Ni����	e"H ���L�}�������'��V:�R\�v�B�V8��H�\�M0;�X��B�Е�1 �)�۞��:)7A�@Gr����K��
oe�okQ x�%>G7���-tM��ˇlh��j��S�X`͛���k{W�f�}���h\{!��f�j�tB������������(��h/��>nAO�� ~�&`��[J#	c�l�Z	�OH~��	���N��K��R8����v^���3���)B�)(����nT�	q���-1�38�G@�$�vL�>Ѕ�\6�#��&�ӋP�L�j��s� R��p� �Q�,f�8�z�H�m��j&�2��U��r�ռ�*�0�|�$,iq�e�rCW���d� �� �9�?���OOE#;�1��D��WwJ��n�V� ��~����mX�Qy�1&6Bߑ?k5dӝOůz�H>}*Ժ}�	�x��=��[�1��2_!�HJQ����3��hY��\8|4�Nzt)#v��5���Ȓ����}�rY"Ú4�L�VziIB�M�ZNG���~QjQ�� �����Ե�fkއX�56�Vk�$I��$b�\BZ9'�Z_�*���+V��3�}���}���b��y����䠌c��	�75Xw}��!{�ڏ�Ho:����5*�7��,�K���0b�&��2+z�2�Ug7�߾E~+��H�Z��4;Mj��"�^WO<(S=x�
3��A1���N��o��ǟ/��$	��Wؙ`�٥.a�7���3�[�sjN`�\�|�é�TY0�'HĒ�nYW�����&��9K��&7�6�",�qA7b[��Q����)'�9b�/�����qUv\�� �{�iu�̢���<]���-����9,h��_"�OA.Q(�b{�*^8���>H���������q��eI&]��"���p,2S��Ep|ݹ�f?m�du�����|����}$x��Z��c���D9:�����p ��S��*m����9���F�x��?@����<3�{��D��ЁRw�I��ݵ�)�j�5�6�6��zn��`t�z�Boǭ͎zAQ�H�+�状��O��K�4qO�K��"R��'��o9�� `n���`��Ў�b�mE:TҦ�k^͌j���3��t+4� K�b�B+�����8+y�����g�}�Uz�C1|�F0+pY��(�^k�k<9���r���2���Xg�o�:T�9�	���qC�+"�,�f���5O5	�n�hCW\��f��v�V^�z�H8�	.�#>m �����i�jT&ZhP4p�qL���L��e�b�o9n�+��@fg��_����q��Pl���[PT�0D-}Ab%�_�;�}��ݍ��8hN-�i���7P�2�LhP�h��}1�E��c�����P ����\=wA��,���Xj�����&;�����F������9	\�Q����ZJm����@S=��D�/�{K�G� ��&.\�ls�i�[�q�"8�6Ԫl�a��������Ɗ�⯁��RTR�K�Aӈ�c(o�s�ar�&q� ����  ;(���oD�� H�8�7	��V13�g O������:���u�����t%��ft�a		�׻�a��?�8�G������eݴ�EE
C���)PQ�XW㳮��9���:H���(���lf��r��M�T�x�\P�,uxu����r��GA�Lb��_��A�8��� -ë�n�+��Mr��� �~�P��{��9�ė�϶�J�� ��6N(��f@�c/[�N?\*V��Q-X�|��d|w9��ҌX��R)pv|��q�-�h`�ϪӲ�b��_�
�?��9t�7�C��5��+]��� 5�,o,/�^�&�HI��#,�w������L�t	��߈ģ�w,�n�It��k"��n{��:nM�J/#7����JIC�4o3'�Ej�����֋��v�dGAĚ�r�Zs���
K�)�_Q��4��X
CA��)X�
~fG���&Q��t625�vl��Ԁ�BvE7�3#��.4�/]��F��Y
*�U�ꞝ�7���ҢrzͷɤE�:l�Y>�K��}V��U�-��s7�y�K[�4ʤk f�W��߃P�����}
���=ǾD��N�O�0�8��b9�4F.��s,��a����@��v�����zP$*�m�Z�/�WX��lsk9���<���$S�o���t_7�ۆ�Pq�����]==�������-_D�4^�lv�Eu�o,Ï[�׉��c�a����^������I�YqSvX3�\�>��	?��-���I��0�ln0�u���3hG�Q,D��p�gя��L���S��q'5�)z�RHC���������.Ɖ�1��)ե�@����&t7Q�ȳk^�k�x���>.j��J�/��f~.z�1N�$�,�<c鼠�Q(�hKH�&m8,�T1:�b�C��P�� ��<��t���g������'���J*���\  �h��
!��Q�.�G��nΑT[��9*bU���KG+Q�'���N^;F��i��.��PI�᪢ZU�9�Iթ��Ф�1,S�z���ah����${cI�hD¤���������&�WI�v�sݴ��ӯ�3i_��jc�MA�b�w����t���6�x18�>����+���LF��'w�U6T��/PU�v��/��c�(�3�ݬA9�[��4�V��;�-���aXH��Q�3��,�B�(�q*�g/������Iu.Z��g��A�aa�����<�'��sz6�Ԥ�z�e=��	��v���Ju+�ƮW�9A�k�a�$�f��?�& T;��� �A́���ڷDk�/4.��Y�A��2@	/[EG�8�2�<.���`[��?:���|�%$�tc�0k4�X4{ ��~꿑������t��u-�y��l�{�pf��Z��4�Þ�w}��U��_�ϝrt�u��!�h~V�g��;�EiBxT 	���RUɣ�p���d]�̝|�X���ě�n�r��$�,V�V�=jApWl�Y�jV&ƨ��[G۪	F)�#acњ㚯=u�.�ׁN7�cb�7�YA�gz�*}u_�3-�h�bx:�t�O���U`��ۆ�N��y�}B$Cbj����/Q�Hg��"}�P����%Q3¤�^XpiG\�Z�L��[A�O{�a�������UF'4�3)r9'��>�0���񗬮�M��ǚ�f�8q���L��?Ē~ֿ����T��xNвJ�<��f@Tu��+\�5Ϩ�4���%��ţ��5�֟݃�}x �6xY�Ǉ��P|k�������j�w�I�d��9�b���D�b�|{���y#Ă	9X����N�&6�����Hz"O��y~!�Q�Ћ�c����L=gp��AҪx8%|�p�{*jI��A����#�d��W���ː�,	m��*C��;.k ��N�BőG�w�|1���^�	|��r�S���/r���[�����߇ <ͤ��^6}�aCZ�I"� ��RЗ��'��l���z�l�0��S�
%^�Y64�$�k/��70�
�����/v�6����$��?<Lj��LQPh�V���٩A��N0�ro�G�����|r9�m��Z�� �=��/T�eHi�E2�A,Z��f0L�#o�Cw~zx"V��S�]/�~��b��h����k]v]�:7�m4���zc�T�b�|�$v1c���y��Yw�3��w|����5pw������Bg����kY=�u#Ѷ�O%ou��\�=����|�D��c �Ё��"T�b�hb56R��~�Ǵ��L=��5�T9Rr��W��H;R)AX�qL
��G;m�0�(9;T$�7Q�o��徣t�f3���$���. X,}�K�Tɞ�Aw&��d������|�i�w*17�𧴐�<��Gz9��&Aː��y*�Cq�!���>������d��oj�};U���<d���S/9��OQL]��n}_;>��E�&{ݳ�c����z�6Gv0� ��\�Rd�K�^����y�KE�����0	���^�$Yv�0�ͥ��Ѵ�nGim'�I^5 �(,ql_I�}H�&3J�mxg޾èٹ�$ 0�����F-ȴa��g��d�]�ѼV�5��Rᣦ�{��$�L�>��\��H}������}�RJ6$�}@��μ��7$��N���Q����1p�f����7L0��S��{љ25�o�L���a,�J��~hM�	�	M�F�V��>ɱ��J�Y5q#����2?m�2���{��న��iZ|�3Vu����w1�;@;)˖ bs3���t���I�� ��j�$f��&���q������AvD_�j�OOO<��D�_��d?��U�h����p����[*�)�L_��+��fhRG_|C�N�����nk/�kYU�-_&
Z���C稦˽Ԉ �ߜ��+���?n��.M���w��yp��Ԗ+nsvA�q���<�"e����}�|Q��P0iͩ�R8l�������P&��!�1�џ�)�jͶG� >0�}�vWOe[�#�H8g���T���L��}/`W3�yH]�����=��x��#���!fe������U�+~�9O���Z����/)���]�^��C�wO�3�İ�Q���c�ΡΉ"[��c��:#�;�Ɂ�=N��s��[1�����e�bQ��:mo^#5�U{@��&��$ ~��zP��r1Z��P,0�a"8A䣝�Ŵ�[�E���),�IXD
����=�j��X���T�
���Rr���},`�=��]�vmo�Ҝgc�(��qwZ��4ی��{����L*F�Ԁ!����O��&�y�� �c�;����0����KG���:�HN�R�?:1G@xx�۫�'^�,wV<���Uc5��ai��w
��m��zO�Xc* ��{&2ڃ�I |�1��n <ٙ�ݣ)KQOX����ks�Z"~������2ȗ��IT��R���MF�H�l�d�}A!���``8��/��|��>b�WK�U-�XaǦ���c��u�2�|�j¾:.��b����Z�q~�&A�P��:k��D��Ֆ��{��Xc�����X����}$ݐ���?|�c����I���r�MU@�5ݦ�ٯ��U2��i�L�fwt�Y���J�v}�PD�j]���-�5�P4��G��o��ԿOM����z`M��k�K�5ٶ�4#�^"$��7���:E���F����;d�Xs���/�>��ui���a,��v,���zx|Z�7L����\���9L"����j�� �ۙ���:b��g	Q9��VcM��3m��Yt~78. ��51s��P�(J3Ɉ�:Vo��>�w��i��ĕ���߄�"��I�=���p8,��b&
��ߞ+���~���F$��V���SY]�jZ�]�dS�R�%�&��m|rE��y����cܮ/�ϯ\p�n��� r�
�@����L<�"�xU�x�KJ#u��uj0��"8�!c��a\�>!�t�*(-goʟ����4��M��r>�I�/�e'蟧d"�{yG!!Z]����$|��O��N���1_;�� �c��7V��w�3����0b7�J��j�څ�WA'm�G��\*L�'����ly��6q�oNք|le�{֎�<{�CCj �LP�&r��P�ͨ�>k�M�c��n���?tRK=n��;�p��W����P�~��x�/$Ǳ8Ŕ"x>?*�b�� �7*���n�ߵ�M��[��-�L�?�z
+ɮ鉽�$ <"���f�=jO+����2���<�������.�	R7���do+�է���.�b�A�g��s +�/�C.�� λ�k��P��r�4A�W׽��>uG����l�����;���l��s��Sf����Er�ǉ�=���**����.�g_��a��G�Ǩ_�ȋ̦�4_�,�b�:CgPi^[��r�="7^ws����!�H+X����;L�J��,�2�ڒ�|��
�QY��Gj��^z�П�i�'�hKʆ��y�f1�&�66��� �hv�p�'T�ha�QX5T���y|�0�)8e��"7ɥ�8oG2p��;\�����‎{;M�ľl�����[x�[#�D_z�w���R����UP��� ����ܣ��^����<�4�����\af(j2��/+��R�Ex����ʦ��A���z���}�&Pů�ٯ��v��������z x*�q������tA��g�^�+G����͍{�[��kN��nԷ�~��S�1��:>]+W�Zi�\��8L�e#�F�hYઃ��*C^!;܁o�|]d�t��/������#d���z�U�'I$�)�N��.V���`��Ԯ�KW~写����M���L�Z>�V�o�
3MX4Jr�:�l{�4H6�����e+b�T��rdݯ%�:s�lAu[��r�=k��_�TQ�g3��Q�fo,�PxD�;z�t��	F([L9������Z����͚0TD�%��C�Q^�[{$��f�6��.��8��X��yx��\���r��3Z�[��-�ȡ�//��ܸX�J���������<4�4{g�{�O���\>5,��9����[!�ғ������{N%�J������j��f�n.�yַ��~H\?X�l��KO3���nl$㾋��c2jo]f�"�ru�e+ܓo܅.3�֧�@-��ǶO��DЬ3�n0�4�dĐ��"��C$�=^�ySr.����-RJu�o�Z��Lo2H����|jrnŶxI�I���B:��;�9�0³�R&���w$�� ��>������p���7�H����?��5&��� ��C�Oi|�5�m��r�=�.����/���@����x��@9T�� ��X=Q���(�[c)1J�H�[bn�/ƣb1 b4�u 4�?�iʹ�t��Ÿq���G�xV�j���W�d�iSl���K$iYe�~��O�"?�9��OF8��.��[����L�~�a�D)ˀ?�� �&�@���^��cI�N��@S���T��O�C�seJ.�m���z�-��,�.��
T�z�-\�����I_���k��%JZ�@�������e,n'�_����!����1�c�N�����0}�Z:]�8�9s��̳w�e���1Ѵ4�#����T8" ��J��2�:@_����A��^�`��X��iK�өa���>�BV0TM,���t*�JH�FYZu�c��_
����U/ɥ����G�vUA(�f��b2�:j�Q>�s8c���t�3͜~_of3�?-�Rۏ�ҍD�����_(!�~,�.�����'fR}��)�=���9�ø��p��?��*���p�H/k�R����X�p�ӓ?c١���Xe�7��i���>�h��d��*_V�"�*�rc��|���D�!��zNl<�eb����N�����OH�NxէT�n�ba+��M��Uϡz��3ۨ??����等�_Š�(y��Z�J�K�4���+��}�@�bH�^$r�J��;[p����W?���D�V�/-t��s4[W�n����$��`�UD磴!
6I�x�2�?���|P���M�DT�^l��P�f�����B���s���I��,�54���w�0����O�y�4��q�(�?�zSc��կvW:a������8���x�mt<��+C�0��������Vj��J�WRk ��Rk�Nǳ*�����w�I�°�����j�����fN#�R���%al#%+vͫHҾ�w�,r-	�4U�����Ż$"� 欲g[!=������	E�h.��6xj�G�C'��l�X�`	X��n`֊����*�S񊕿�RTl�f�����-Ľ����~
j�έ�w�m�����H���CC�����H|7�2{�*�[.�\�B�WՊ b�]]3�7x%M�yۻ��Y�����w�s������ౢ�a�� �(�f	�ϛ�φr�6��x���a1�s�2un��~a�o���Xj�n[��E�I�~��0�/�P$��"�u�d�YH��̩��!�Y~{{��N25s1�WԶ����ln�k��ɼ�M��@K�S�S+��f�(��ÑXo�)?=?�W��d߲G���7)�C^ZϷ�f#ņ"x�Eن�)��܏�����@��ko��0:F,N1�*���-u�Q̞�Z�d�Py༳@���YA0�N��U�Z��p8?�����L��]��f
s��H	ET�sS53[SP��:��b�W $#��?�µ������ِ��6��"�J��|0�����w�^'�<]]��nSz��"���g|C�fO��V�5���}�{�߫��oi�
�O ��q�X�"+wF�I~ In�	��<�/"���u#$k�b�X����[1g|lQx
�T�#���leo���1]�L�7�p�����E7�����eh�K�
^-�4��k��yf��;Y}?�x�gd��I"���sAXf�j6�R�4(�����Ms$�a�nkg���P�f�����y2CyT�k9�6/hv4� O7o_��v䛳�_�	$C��sQF��QʢĚU���T��*6�ty�K潺&6���Q���vx
;pX6�̦}�����s���'������D�S�ox����Z����RJ]��s��n��Ǎ\��<;I���w����
\�Pq�lF�5:�xS�|��Ǥ�A�nU��=����C��ߵIPA�.5S�M%4{{�̟���#_���B����k1_�cCEt�.����R�K�8æ��g%�fս%>
�{���v�6T�T��@TO��P�h�	�	���h!ğw��3��� ��g���Y<��f��d�y,���:�WF<C$#~l᩷�k8��i,����?"4�Q؂�\ݼ�u���a������q)\��8$1���)<W��������������M�Y!��H@�)d��������#r�kЯ�-�^S�{x`��wQpq�x�,�n��Q��+�
 /N�Y���l.D�Q�6�4�s�C�/���&a�}�>-D�m]�]������G?&j��z<��]�5�v�)��[��F\�G���a��ػя����$[�?�YoK�u[V̻̾�L4���Kul���^i�(�՛E�����^��a�W���W*��p��C��)?bX	ߕ"q݅�:W��øV�����5/U���b,$8�V��m`Ώ�\vtΒ���΄�������{ї��Ob�O���5ʧ��U:l��=1�v#{���7�#���>ʄ���?�d�E=���h�(}�j�װM��~G��߅vd7�><­#r�J&����n�s����;fx!�bJ%��A�_�����P|�&b��p�>2�iu�m�븐�YK$�!l��XL1R�#n1�%�D���W�JF� 
�9��a����&�8�V;JtE��.�x����Vc�B����6�ƀ��A��N{#�6q���w<�`�6�-Y���� Ҫ�S_.�̓yX(��y|.�L{�&�1�}�Ϙ8�z�u��,Tc�G=t|��x��?(*<B��_J�{y���JA�o����!�(>�o�����^�Ń�d��}^�z ����{r��^�#�s��y*�c����!A����g�{���U��E��}��sA^p���+�i�w�$��/�oHno���Kg�r&��n��y��������q8�*yyX#�Ш��.G)>�/���G$J}ZU^���
t���dQd�o/�>��׋ԕ�u�tϲ�F'���s�!�(�T`��{򎛟�@Ữy�n2�w�� 9�GY&���Oč���6n�-A%��{[��k����Or�L��6bi�K��NP�>(i�=�eH�Q ��'�J�q��E`�;��pc�Jԣ�䟆�H��;L�ӎe�w�2S��wP�#�^�E�d=�2 �^���>�= {vC)1���Ÿn��z�����n �5���N_0�4���T��7�QCn��,�]���F�F1&����8Ç�8�FMn����2#%5�o?n�î���/5��K)R�T��)��m�������o���Zq{Ԫ�ٗ��hd�/bf���5��ԯ�����9�mJ�P��ir�|}�O��<�n�>��;2�{������1jԏ~�Zqb:��m��l�묃]�ϛ ��nD�ԲQ���1�2Y��Z��+��`��`܂2��a~��4:H}��W�c��jF�L�:���ݩ�à.��]�]$�G��A�Y��|:�� ����믈�*f�8�?��X�{r�7_''�� �ѣ[L�`A���I��(��fU�����l���ט~��a2@�~��KzDp�im8[��q�§��{���0��>0r��`�v?�����A�����c��(PҖ��;�kغ�ik�
����#��B�h�"@R�Z-�p�!�W�͌�bu,Fy:�i��$`0
�X���3+�q�A&l��M���|��e��/qO��ŝnmJr���I�N�|b���i��5PY?-�w	].@AB����Ԧ��r�AB�����ć-Ǟ�\Vפ�x���sq�3�i�Μ�"NOף�*y+�|�~Wy��*|�6.e���*�aA�I�+�IØXG^U�J���7��I����î���'o��A��8�5M�)B�hT@R-EB!��Ɇ�G�;�	��qF�CF(��O��]J���l���3󂕵����-�x3qz��4.�y�si?W��qF�Lo�}��7"�0����	�k���k�ٸ?fGyď�'�'�xk���"��#r����[Fp�������q���̐�`eݵ���y?EJn�~�9f��S�	IJ�W�mM�e�����_	v*i 2o�W ����l`�M������7-��$wo�ǎx��A˅�o?���[��1���uf��-�6)&чW���0�l98d��J�A���j�<��/�ք�`��q��6�V�a��biS���J��T7V���:_��L���S)�vg��AD�&�e�[�:"#6}-���)v�^>wa����L��$8�F��@��p�2�i������r"-�u��k�(��Ug�gPUk1�ޘ𒲿�����LW���$�d�2�`�:��b�{��3���Ư��ha�櫒�a��!�뙜�e�۫*Wsݣ7�dkf!�]}��=r��-Paq3V���;��쫤��0�DT��i�>�f�Fk��^�d�
�Q�ɼ��v����c��[_c�I���4�.��p%BF��^2�I�������oo�9�Z��_�ݼxd��5&�V�Li��/�>����zګgäQ����T�)�I���7M����nD�R��_�r���w�  �7��L���\�L�5<�y��;��=�X���,�($O�������V��c����W k� ����gkaߎ��_�VX���)��V�L?�#��&k��"d+�1$wEK>���+R�yԫLkN�V	�7����3��a-/�2ɚ�P�N��;�������<��͗�ʃ��}�Q���=<�Bu˦k�}�3��,��=��U~���QA�=��J�~�4%�ʡ�u.<�v~~7���J&о�7��}Y7����}�x �p�gծ&��F\c03�Qo����ػ����Hz7�1� 5 ����;���͌;ƏY�	v���o-�K�ī��Ik�|�*a0��B_�`��B1̓J�k��5	��,/N��	���-{3as�%�:�C
�b���ax��%���d�ڗ�P���1��FLw}���fu���봷f���)���)�>ဇ�_u�!�����	�k����\��8�_1(.�T��.=�㡦ZUH@�S���K���g�O�b���	�a��喀�Տ0�*L(e���L�q���A�HV�hj�0�B�#�^�.�r��n��;(�
��1wZ�|La{ũ��I>��&��?E5]��)�-���l�5^!?kU$���ݫq4�*$5 �'~1r�v����Ӂ�) Y�_��~�#xW�c�����Uxi^��cm�k���&�$0�u�/�����E�>�4��۷yx&��'J���%z3�7���'6���=������>W�o���Yc����fÒ)9?�[�<�nM�"zn����Ag��"<ϙs�hw�͉wA���Z~�� ���y��{�0'���V�P�0>%*�6�13�:Y���ꡯ�v��z�F�1&|�'t��� �U�:�+�#���6�T�ݡa�on�p�}��qEW4���)�eHlׯo=���}�C%�s�&�ΜJ�1�8K$Ypz��p�2kVu^"y�-(僡Zv\,��v	�2^P/�!��-r��1�I��
�R�BC$)����{U��;ֵ����ݜ�	}6����^�����T�?y)@c�݆�����±u��<��TSlBw�-l{(������gV��� ���[����Xc���v'���V�4�o, )���TS�����j���1˛��H��N�(�.4�����N�t�w�-�E(t%�}:����[���
+;�ً��\L{|�7�y�kŗ�/M�X����No��A$�Iى����S�ȘS�=,e���Ӕ�7/r�'�B�A�Kq)sc�|{��zDJxq��x��:Í�/����B#"fҳ><�����nC��atg��D�=F�zdP���3�@|�YY��l��L���O�ڈ3~�'��1R��,,���#����'B)2{�(=�f��HY�}� j��6'L��S����}T�ax�^�DA�җ�N�t�'g򶷲1eS-��9�Q"�nA�c��:p��]-t��3���<���ǖ�&����SO��ꯄ���Y�COI�A�F%�b���<��sB/��^-.2����W�dڤDC;��vc �:��K��)����~.V�a��i	"�F�)a��{ =�t�-�r�-���oP��e*_�^	������T�.�uӗI��H���z���3������(���а�q�rZٷ�Q����#��<:��+�U��.��a	Ry��b�
�%8�n>�I�cJ�3M�mн%�]E���{r������R:	��0N��Z��F`�*��P�۟+£�:2��N�`�b�ڳwfI�7�&_��e�G� �hQf�#���A�g/��O�!�X�}�'���wp��=�D�����R���>И�,ǫ��o�05>�T��TTY�����͉���eD�0��ۛw��\ܰ���Ԯ g��[ǃ�ı��L����}�fT��_ �;^L'h�[(��3�с)�g�0�)�,��������J�P¿'cs��)p��NDa��f��_1h�+4*�T$(�e�y��$���SQc�ʔ�ɵLN�j)�׮��J9��iT��a�抈�/�Oc��bD�t��;j���l�u���SV*y[3�0q�Z+��M��O��	w&�4I"g��=4j�p�v��ҷY2��+�Т�!��b�A�E��'��{�nj� BΞ�����ҩ-tTa�Pޘ\��-�q����.R�����0�M$��#�DX�+�/B-�Xn�7��nyJ�����6h��4�)a\" �.`P��b�>���!�����8�d�˲o�^&Q�u����oXSƟp
����̶���t��NVN�@��M}��lw�:[��O�sa���q�m�~>����O�^ujYU�&3��<���Ѿ�4$8w3'�����l�}t�[0�����E�x�J�����#�"O��] /6��U�kB�j��r��=�	���X�+��]�ZP�K�4	q�ܸ��6hr������G��T�A�T��	KP��W̺j���o�����L
��11�X�D�[�tϣ�2�i��gW7 �����'G�8�datĴj��D´�c}��uQf�ֽ/�bq�Ha0�)s����R���x"�pT�	V
�˛��,h���
m�U�m+[��dS��A�x��G+b�8}f%��M�]\L۷�$�7J���Sln]mh�:z�s3��\f�+�Y�-��1p~؂ɘ���o�P݄7ז,B\6Y��/�*�=�����M��/�}
�5��MH<�H��2v������4�^܀w���N�J�ښ�%7S�@����/�p�(6�zeDy�_@4�swC�WIEc��C�.^�zZU]�B�Q�.+��^ 1���W}�{������#�8+N'�6n�:l���>�tw�;���o��7��C�[�^�rh�wD��O]���VrtvU����;!����g�{煊��)�8P3�u����eU��/�k���}���E��ndG�;f�yPI�]�$2G,�b�8�r^��xle��ݘ#�3єu���1�_�v'S����. ?h[��6��N:�
5ua����|�����&j��:��D��ph���&7Hܭ1� =bC��jϢp$��DK�>^U�3���ÞYey��H	��>I��~0{����o�x`�a�5�\�̂�>�a�_Нt��w�K� �MK���H�r�������x6]k'I��PHJ�gy��2��nk�q}�G��80ʼ�n {���L=�Z���֊�_��� ,erA3��3��Ҟlt�sO���`�@{&�f��u�p���	C�74᠄�-��+�6����Y�Z*mGUZ�dn��F.7��$2����X�oz��:�-��6��Aޠ����o^������d��2h�Y��Q��+ԿZ����%6�~H�8�� H�GM�l�)k���Qb�E`�Kۈ���K���R��-�5�����lC2eeC�J�̿�l1jpx�h,Q��<6&�mʤEj���mEH�&˸�����p�M���wT���=jJf	#�%�Y]��;8=�O�	�|4;c�6Uw�a���:Œ���\~'=��)�ڬ=��%#��M?�G��÷��DV�,�Xq4�
�����<��@�e�����wY���Q#����JgI�Lc�=��͝;��ٯ`�L��\����TP']���hh���z���s�쉲�HP��%�C}����tx��T�����2omWm���E����D�9)}d����Y������
3����9ݺ�> �?s��圃x�\vG=�j�j�x1�yJ�o�8������~�*�KN<���~�ن*H- �6[�~�Kq��,%Dx��p����N4�`M�0/ɍ�"��!����4s��ʅ�� �ڐe�5�sЖ�����p���w��zWmΦ��M�5��)d7�v7`��ED���*���Q�_����Zϻ�/vr~�1
��=;����K�c�ֱ��>3z�jv�T�i�q��AA-}�/"P�*-�tEK���,kD'?жG����-T��s;�2���k(��'ƒ.+�%ةJ�k��P�U�^�0x!��A� �êӺe�~��sl�D��!����â�?r9���vM�5��{���4�_ӥ,�Y�C�OQ�n���}x<z���o�Nu���.�	����D��Ҵ�'Qj؄��Ό��'�C��)�9}뺮!h=���ѷ8A)�y��n릮R�A�9VP���DM��:��[-�>�躺�S� �9���i9�+�=�p�i!A$��r>��a�k��a�I���}iв�s�Ёd��|�p�����e9.fQga:\��uCn�3098�Iԓ
���x���焪t�l�Y2q�@ &�>�<�2�~�0z��$���U���-�>�I�:&-�q؃�1۶��K숥�ͥ~R����2�h�7yʁnb�`oЁ��َ���m��N��$�Sx)٠nY� [�Ȳ�����J��� Ǥ֜�(˩A���0fs\[��!&GEKG"7I�=yO�j8���r�t�#���ֆ����_�?���)�1��\{�&i�����C���ޘ,G�T�b�1_�N��+S���d�Pچ7h1�Ʒ��#l��K��'���rOB�-]"j
��� z�t	��E75&b�nEFG�ū��Eu�p�s6Z%{�m�Yc-��Qf:	޳���B��S �b�rm�s@`~�!�h��ծ8a�%�?G��'R�߾ s����� W97Л���D�N�)1������sۻx��C}&������X+�Z�w���gc+h�Ǌ����x���Ȓ�����zH4<A4�e�~Mݛ4�j��&�S�d�'�I�ᶮ��e�0;����	ܲ�|���4���FB�O���|JP|F��H�ىB��`�r�!
���(~�����羜cSWA�Ԛe�/!�[D��/y��h��,z����
N5-�-�Bj�R�{?�|$�m�}��k/7���]rKm{�N��-!y�w�[V��k�_�Z�b�G�N$�r��ځ���r����Rڢ xpv��-�T-��������%�°��-�ف�����i!(����s;��W@������eh�����"�e{ q��g(ʬ'2�e�֣S��0�aD�7`��V@�6ʦ�� �r,l�ժ��8���d�c���Va�(�f��~L�<�h5��]J�/�?��	�o��<��x���%�޽�M�2�O%tկz�w`{/����M�b���������� ���S�;����Xe������T�#~��|�aT����%���qS�!)�Cp(��M2��n�}Tת�ؕ��w��P���G�'�M�i�X:��K-�~��m-I��#3�u�6CBFW�
��Q�c�q��EQH8���j�x >]���+b�9�Imr��$x�M����j,_Ԡ�J�#ۭ���=(i���Y��)�%6g ���xg+(����%iHZ\س�����d[%}�s��S�|�3lm"�6��b=��'<l�W��s�<0���w�\~�[��C+�������hU�@4W[]s���Y�`	4T�4�L�O"P�2?�XO�ls�ܲ�D���º������"��ʠ�}�|�v�"	Ng������jD��0��4::�{�~x������A�x����18�&��4�G�6"�֔���´s,>����c�`�z�l8'Xo�x�{ރ.�΂ ��;��_8�@���4r��&_���.6�
��8O�x�f�sP_*\��ڣQj't� �����w��������s��L'��p��#�6�f4(�T]�i��Vg�+�p��$������.u�p�8ˋp_(�%N#P��6����J�p�\>*��� ���7r�ҋbT�7�]�g��$��{��S�� �,�=����z0����+�.�X94L�|���VO����� ���^�<
D0��-+j�!h.s�+�\z�[��#��|<Mm�jVԴq�׀3nR�r���| ��?�Q�7�k%��[A<r�%�Dh��M߰cu)FD�]���uIa���1H)g�_���2�M_��$���xa�T�F��kJoD��Pq��޳��M�ed4�+붔"����N�\��w��D���a$��~��Q���_���	��ٌ��V���.�9���٭��n�������zsm�����1��3����$�oAk���;�?��<Bx7.���S����4���aOks��"����P����(O���ڰ@d%�j��ϒp=�Ԍ���F�b'ñ��p�Cm��X�-˖kNPe����	�u,�&
���޲�P�fg�M̀{������DO�������3�6�Z��W;N�@�o=B��K(�`tԣ��S��L^x���L8�Ci,hK�&q������	\+Uc�eo!Q\�V�1UM�m��<Nƅg�_�	�<}�2��`!�x����VD��7�,�T�*�la��"��΁��rU9�|���X�.�����k�iPL9��7A�jŌ�E�s�bׁ�&cj[��Oߔ
m68!]%w{!��LDj��)�}����OÓJ�b
���vm���G�NＱ����	12Ο	Y����a�Vy���Ͷ��A{��`F�Q�{�!%�u��t u��?n����d������"{'�<`���J�킃[��$T)�R6e�7+[�8��0�
� R��q��Y?�&9KB�Nz���6�Ϊ���D��^�=N�ͷ2��y��)�x�����SEST�v'��;����2�%훑C{�^@�E�d&��o�5��8̚�I�19�Mޮ���Yfe_��䴧v]&����?<Eaya��b�@�<𕻍�	d+Z����S�F�^�o�I��x�)kI2َE+[���ǤI�/ݐ�IP�(�y�m�z�`K}ؗǢV$ك϶(Ҿ�oyu�S��� .�+�C2Xrų5]��[�B�0��-3v3d�m��_�^��v|����e���� ~[�Wu�\9NH�kSi�n�| z���@}�U��tB�r�<`�9[6i(�x�b�]��ܞ˲����9����ómK���"�zΑ8@�S�R��t����$V`�ce����*q�-��Z�B5�L�O��YcJD(H|����%�Q�K���������p%5{ �����]\X1k��Ζ��ѹ��:�ᮦ&��9l�S��bZ<	HF(�J��d�-u(58���,�������7�ſ��%8�b��)1�rD}W]#��LT��g�0�_7tK�bZQ�y�ש&ϼǌ�E=�}����m4v6��5ݒ|���~<h��Y�0X�+���2�R�0f��	�i'�8�X����x��<#O�+<!U�q�<��y�݁�Q��m\
VĊ����s£��M���D+�c�S,<+m����nh��=�Q�1`C+��C��$ ^e3Z'��R�͟��s�T����6�������	ay[�tz��dD��^�5?-6���>N���@0�4?@�pA_Kf,�-�yN;�*ʒ��ѬI6� h]��� �|�Yf�~�|d�$HXtF_�h$�9%�B�e���= �	MQ�PyB�LRy!Y*�{VYt�]$�Ā�lde@{#٨��λs����[�		��s~M^�K��bt_||ٸ>z*��A�G�)G��}��#���!Φ��]��33�p*Je����B��t�dXb� MQa�^S��t�z���ʁ�qV6�p����V��qL1����՗�rTw�"|d8�
:��~6d]h���ϐB��Z@�ۈkAN��<�l�b�C^��r��>Zy�:�;d�E����m�c\zB_q�s�4�|2�b�Xe�����e����n�w*[3�.jـ�6�6��#�����Ʈ1��7��/P�1�����!�m���G�qB�ߎ�д,F@�_������U�-B'xb�X-�� �W�\�:7@��G�)��m(]
E�o���| o��.Fǁ.:�(�m��x<,�5kB!p����1���#M1l�x�myK��fq������"�dojU�|
��	���U�sY,�l ^�_v�}>";���-��-�:эU0�e�XHsx9?���kl>;�<�i���,��҉��<�2�[Y~���Ѩ3�<��=��b�X��x]��ǧ���*��uȯ�_�W�N��zCxE��'��/EsdN�w��*�^X�]n%Y�Q�B�l!�f�%���߽�wv�.Qə�9�?�a��P���FF�ǲ��~	yȼL	����|��10\:]�?�w]FN��"�^�#N���Ȣ*��(8nөj��p�JR1Ay�W<����	�GŽS������p7H�}�b0��}#��~Jk�*E�5�Ϯ?V}�F���\� ������ d���n?�&�69��"v��Z]��4�7���,2z��NwbF�=ի�6�6�K?��T���*��Jp�-��KS���q)W8x1~����f�h�>��JQAL{^��\x`�P�hU�L�H�w�H��lܣA�7��9ۏ*�Qj�t��� ��L&VJC%jwmW?�>�������?2�����s�N�Ʈ���_	�f]b�O���d$l���AU���o|\���\Xl/�__s��Ca��X�k��큨tq E]�~�a�r�i�r����E�����X��lw��DI ��¼�� ķ���x��!�W������c*�aV��s�I�1T����I.a��V�B]Pq�f"-��K��ݥ�~ֹ���t��i4��ׇ��-3"���;٭1��Zg2NmiW��9_�Y^�)v�n´�l�/\�Gj�op��9#2�7�I��uQ���g]}�g���N��F�X�X߃ֹ8�t�W�0������@S���SXcx��4�z� 62wɿ�Sb �ů�|�j�9�@!r0*�R.>���[$�