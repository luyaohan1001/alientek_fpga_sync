��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ�����D�!Q�*�>d#��ڥ�*Q#���ߘ�S'�8k�H�����[��LX}��IC)�4��g���lh�;\��<<2�Q���5��`4Z@��$3Sf	+���c����͝��)b��AM2iL�,�e�>Q���oU�kd�Q	>�R��q�������������%���<����À�m�x-*`�uiÍM�5�s0s�h��!5����͟{�g`c�y�lHlE�D���˿������0�JP���J�R���1>�*��P6��lpF@���N��)�bq����=h׃�M���\ש[V�����ꏒ�ʪS�U�@��O�(��	�wv���M%B6L�җ��si�W����]�+���pR�}�[���!ͺ0���[��=>�ΐ���'�U�U�b���ӗI+\dT��s��(��w�X�Rs����Ñ&�֙AB�XQ�'�� �$�W���n�0YAcY/�=@��|���0%��?�M���Rp�hl�r�2�
8�#��V���+��驹�3B��ϰ��}�8M��3_�*�°s��=\D��j([��_O��d��c��V)?�y�)H�>ɜK�i�m���7|���	}8��q�|_��7����8����냧��A��}h(��T�{ �
d���^:�a��x�,�+��xώC_&���i�o�`��h���6
�E�J�@0�Yvh�����&L:e�0WR��[�&)z�m���j�e�6�;��c��qia�g]�E��W5O����SG2sohw�S�Q��`�{u1�)���NZ휈] s㙠�������"���8_|�Ht�TO$�$�\/����2���s��2�:�i�L�����Pf�����&S����8��7Ҩ8����/��XCE"�l��ؘ^3�I{9"�{�&C'}���@H��T��洶�f�����zK9n(�[�����4G��p4�����cx47��K�N7�����}4�NK��ka���������i�=L�On(����-��^��*���=a���z@E���,oF;��XmF�ƀ��G��B�胋�[3K��28�9Unj���iP5�LQ�<�Ƈ;��	�Ð�UC�̖eb�ї@�ӌt{��S�m[P���R�(6�iRm�Bt���zz�ub来�5��AK�����%�{��zU#��28�Cf��"���{�4l�fr�9�P�6X��[��๣삢)�ѽ��:I��*�S���Ksj�e�3R_�EB6�9�j!��j�m' ~Kqf��l��Ss!�Zn�5���v~����'���\�����<Ĵ�֎�}��9��+� �l��kc�a�'�͘~�(��X�/���J���V�Z�6����%�S���<BDK��\S��;��7�du;GG���T�M]R}Bٱ��6�7�n���, $[�h]������ݧO�Ce6���|�8wa���IU�� �ą5��^D�/K�J��
�E%�fض�a��A883�����Ĕ8�SḪ�t�P��R/�\�r�m�B�'�ښ�&P��ɽj2_��fP�4j&�@�v���#. љ�E�g@�a[��@b����/BSz�R�xw�o,}���U�V��	@(�k-%IL��6r�� c��
Ҍ/0�ҼF�֊�lЗ�^�������Q'eI�����O4��*�^�E� �3j��8��4����	xZ�Lg_���$K�`��{����!+v��{tN`RH�������0�X&6~FG*gX[} t�]t����D�������WcA��vt��^P�}ӟAD��>z���Ve ��L:�0x'��@��4C&����H	\׵ښc0<����X�*Z�i�>�S� �]�_c�o���QD1�����5�ힰC]�V��SM�p_�i;_C�ܷ���`iE��6��ɛ��P?> 
���A��Ŗ>Jtz�5�Z-���˔�&^�;�����o d`��{<�5��}b7����T�v��'�w��[m���q�E�J�k� J8��v\$�9�cFm�����:I(4w�~,�b)X��2Pc㬽@g���|�<Ӊ����8��� ڙ�5�����eR�Pr�E�\�}>[#����6���Z@7W3��o�U���
��X֡�b�y�,ߑ�V�=��(y�h`$�?����]���\�1���
�u��bh+�(u?P6��qOX�<�U;���p�\��	�rjs�R���ct��q{0	�2̧�g�C�=7��o�ū��7aBoC5�V_ѕZXS`cyp���Yz5���Gc�}<1y/���J�v�����ƁP?�z_,�
9���V6�[�sM�F�7S��r��t)�4�X����������w���i�������������O���KC}'���յ��}c����G�ܰL^��@���G�Tɟ�I2�%�j߄���z-y���%�3�D݃Pޕ�a
2�%ҍ�S��'P$pn��N�n�����D���1�rw�*�����-^m����8y�!ɥ�nڃ[b�T��(,��L$�Hc�0���4�%�B���^7�����l��*����9�؀LU����lN��O�eki4�CP�QM;��l��t�,s�L�+yA��v��z/��_�iy�0P6��nS��i_,V��d�B�m�آ��q>�w�U�|�껅�`�)�/)��̈́w�
T v<lI,��v��ߗ��L�$?t�R��튩�b��i���;�'B ï�����5tZ���a�	�A��n@n�����8.D�ћ~��M���$ͿvK@���~%�p�)�U��`&�kky��#��]gx����4~���ZV�V{ �w�Wm�OAQ|AO+�ǰ1L��nU�̂�dJ�a�~""�g�3��w��!��^4�X�Ww7���R^�ˬN��Ԃ��W��J��;/v���.z�����"�}R/)�ɑ�!���)���C��^>%9����M�*�>�4�j�����h�.���1�Q��5ڙ���ƴF�
q�M� HN���ގ"��h�T�^�OM!=��(�'�Ⰺ�[`Ŋ�u���	\c��K7\�w��Q������v��|4�W�榋c�cS��}��A��ud��|��J���O�'��N+A�f�n���^Y��8$ا���Sʯ�d��-Y(��鑌C��3w'����1rԯ{��]�|j������ �E�f�l�:�ig%�5�u	� R��9��Җfz�h���-����Ѵ�b���'���b�+��hc��\Х4�s������rK��I��[ǆ�G�pl�A*�����y��#(Ik7�e�����	�o�Ǳ���v?��	�9ǫL�3�]��b;n=��OBOU�t�]pn�Ȝ�w<���O��Q9���T�]���7��L���kJ]�E"P	j��R��S�.���37��D��B��N%5Rk�4�1�D^b�Z�֬O���)�����P�u�oJ�%<��*�A3t��t��bg.���|�A�E��a(�<��Vs�`Pl��I�u_e3�S�'�M�5�?��W!�� ���@�V"�	"=\���՛��{�q��V���*��(_��7���i�g��5�����!�9������ž>��]��g"{\+]Q_�u9��	�u̖��*^yH�~=[�5�ju�$����������d�5��)hB`}<}��8T��0��8B���́P�#=(���*�x�-��g<�����kQ��.���I��%v�i���>�'c��]Ԇ\���/��I�We�i����I��r��!0�DL�H��G
����ޯ�������f�͟q�s�rYs\���QY���L�&v�}YsK=��S�8-���;��o���cv2�,$e�=��cD�Fl���F�`p��d�z���V���?������x��+���9��|�����%	��i�!'O�5���m�6R��.�<�����LBꆐG,;�n8CYt�c��V78K�%�J,�Ö�+�AB?~���,(��T)��f~<�)l��8�Z�k\��t{z�b� Y�K��z�zk~�weLșCuM�Su�����׎e<��E���[�X����K(?�A�Z��_��r�3��c>������MEǱ��������ĩ������A
�ߌ��g��Rǹ��u3�)|sȰtǲ��xg�{ݦ��)�Pʧ�e[x�&=�+ƙ����
�ȋ�om���Z�(�>�����1�_u�B%�j[L�[0�أ�~�,f���Ԥ{Ϟ�ӵM�Gv+/���s�y���Fh�`}*�қ_��N�k�ӛ��`e�O^6��uG]�PC3U�mr��k�k�D��5�%��J�$y~���N�Z�m#|{'���F[��?ڳ�;�����<���q7C�0�}Aя�< ���9��r��y�Q󑗦���� 8>�gfh��m�������L5�H>XO-oq���Uj
�[?T�K0�)�ǥ�0�FFL����sp~C���%e�'�ǒ��f�P��e�޽��O���""���LNm{�bFy�a��ߜ�Z3_���
_�'�ZT�ήt.$ÿ���4��S�:���k%����ɷ��g��-��FE��W�q
��|�]�˻��=Ǽ2�4վ�J�X/�8�g�� ��NqE��Ԭ���>j(F������E���t�;�mF�Wm
�o�x#Do���"�IN�F�*�4p��}�o��VX�����,��_D!,�����?����ܛ�*�X�'��?�qN˯�c�%�r�� �m
]z!�HE�h�o[L�:�{m?:�ɦ��O�lw�;\�Z��dW]��p.~��*���"゘�wI�2�LU�.?}H޸�9�c	�9�b�a)���Jnӕ�=�-� qhq5*�w-��p�d*�KE���l�2$�������T���*�e�p�$�5Ð������9dm�+ �6x��Z�/�[�&��ui����/b# �)��d̰0)�ě�H��ۄ@A�_�J5�4��ĉ�%�y�69\)�����Z�L�ņT��/*EQ����3I�D�����@��I|����'�L'���K�ĸ���FA��_�2ι]t�l~͚�Hd]�~�A$
�"��<f@�����|�]��@g3H�;��&޽dv��d���"��)�u�ۺH��_*�&N-jy�c/��D>iŰ�!T_���z�����&���x(`Fj!9o�1�}��1���/ۍ���n�3���R^���ne��W�r�:�n,�Q$V|���Aa;'�(��J�-h��j��"r�J�F�O�t,�K5B� �=�\_��bm�ﶌ�*��=�>��Nw�2f�\u"L��qy��*ϓه雮���k���udݿ��.���s��֋9\&9*��:���Ա�vz1jG����	���T<���qY��x���=���j�%U����뽱����xj953���+,�u���1�ehe
��ȋ����u�u�f�j�i����nP(��/Q�h�W�힝��']*v �c��PѩKh'��Gߥۡ6��MRq���i3��������N1�9��H����,Lt�X4�@��c�,��'=��q;~`�x34�D`ɠ�ijD0��ϲ����Fg�	�T�$\����#���ZEB�a��J��_ ��݌�ZJ!��@OWF�O~����mHk�����:59��� ���'�����7Z��~���eDȨT��x�ݡ�
4g�t�q2wR�ԑ��{���;};!	�8���\�����F���r�,�Tj$l|k��gڡTgU��$d?�$��\Q�a���¥a:tQg̠_�b�+��q9�ѭ� i���Z��u�h���������'��\�)D����ǾrdymZ჆�˽bZ��: �	{e��rEp�
jbH�j���#�7�I1o��/B�%��lk/�C���'e�U/�+n(|��BX�?w����UE_lj��%ˏ�s�K�q�^A��QxK���$|�ש���tW�6�������A��Wy�BbQr�ȔýTi�z���v���e�"Y���%̨[@�1�>��/�,,%��9��<x"��UԗP/&��N��g&�c�C/�aߜ�ө���/Zk��EP_'��n5���R���tdu��ǱN�&�.;��G��o ��n��y5��ص�<̽��-*t<h��Z)w>D��d�o'�,mÝ�Q3ȣ�L��u�@���>SK�����ܵo��^�&�T|V��T�ZD|�{_MDl�`��,e�R���;��WV%{D��d�sA�wQ��x>�O�,[sVL��{�z�4��F�L[�Aͮ��D޸%���I�O����/"nK�q�ZN$��Yho�P	�Y)b?��$<�?+e)��_���@���	�f`2��s%�|��7\8O̵Gͤ�F���O�4�5������7�a(C�D3���.���N(�,��a{UD��p��<�r7)�SV=XMY��� �`���0���I�K�������E)�lj��³�����~���lW~$�3���s��K�"�zW?֋�`H-ob2�[ѵL�K')�Ƀ5I}�T��3�s{1��/E&~䏔��Ǯ�$�Q�V
N2O��+Q���v@ӐC�vD)f�A<�G[�S���4Tar�2�[%�Ab�s>�)��i�	�8��:_�Y� �[r���N�e7�͜ѣ{a�b�ٝ4Ŕ#� W������b,GW�1��J`���,n�I���TN^��q��k�~�4�� nc8�
������lr�Q����v��5tG�`r�4��VII��VouN�4&g{Ȅ;EӸS	��q��v{4�e�G�v�9'.-Q;]�yV2ʯ��qX���i:[[��Z�@;{�p��S�ͯɻ�]9*�j����n/F��?��������6C����54M{�%j��/�����3TW\��V͞����d��ineh~�lW�����9�M�1�i-��t�~�Јn%������ b�c����@�`�Kӧ؄���A<d	��qԆ5	���y&�ݟ9�B�e߼��s�snH_\DyR�0]$��M~�z�-��S��nn�B0f$>`, q��hg�[7^Q��%Ѳ��g �~�e]@_Ɣ�-�!�5̼�!�3�$�$W8���8�W�!Z�I=h��4ٹ�cdVb�O�����y�*5"��e�j���c<�6���� ^Of�F�)��G�&��K\�����Mn�(6:�e-1��s�VRms��b��8������xw������w������j�t�u>�K�l�G��O�髙����2���q?���RV�;����70�}�U���l��9kZ�q��f�A�ֻz�r�
Ǩ��iynB��Za]�0!�Kx�ۋ;	lP��Fh4;��,�xpR�dq�+�1�E��>q���`.�b,�-���r@�p܋,1.<#�d���'<�u���U*g��I��VH�=��N�J4Q�i���z����U8�d��][�(e���.u�R#��͏Yt��)}j�ż�>>�~{���B�������{5?�]i?��_�"
���\
�q�{	�O����Ϸ�k_��lQ���8c1�	g�]��ȣ!RyB���τ��g}��?��{ToG����M�?Z���JN?fT��}k��<�s/ۖ�U�{����ġ��ĝG1ˋ�R5�^�E�HN&�����P˝�6���e'�ܩ�F�0�q�^"���Y_b�����v��pol��䈓����ҍu~*w	�����o��jT�O���<E]���վ��h�Z(]�,�E��wTP� �aPS�HCK�P<3H�w����;�\ݣNPؕ�Qz�$���b�f���0�Y�/�A��Qb���'��t�,�3����g������z��^��8�n��m��m��3rp���-�v�^�XϾ�k#��otr�:���(�ސ6���`|*�+B�*	>��L'aU.�9ۊ���j������ŋw-A��uQ)SWfCx�}���f��Z����w�����SX�^J�-�,�W�
')��!�ji8m&�����;Wp	�E�0�H�5b#��Ec[���~iI"�=1��;lm+�`��E�J�'�#-�2�u�C����g�WD�L��x��,�O��.�p:$*�&��gi�?��W��;������"Wp��pvYj:�{�8��h��XrHB+}}�7�ߧ���G
HY\ծ���e��\>x����xRB�{�ЪIx�t�sY���Ȫ�ҕ�u2�'~�0i+Ԋ���eYE0~�\�R�`�����	���?�� �3�S�/3aj�>�7tŉ�n_���2�΢4]�T��G�������5S
�?"q����m�ϒL��_���3��9��3��9��Kw!ڑY$��&�h��!��-��&�`-�H������@l�`L���W0�=�V�t���zۗ�7;�O���W�tNWw���LY�P��>�ˋaW6��Ia&%�%���rq��Ŀy_��J�����?���&����v1��v�%��A��w��ݠN�ݷo�}dSAj�s(����Z���o���]1�Ԡ����ս?Sd�$Y1(��Tگ��rm|�'ݜJ�6�@��
������l��E���hSW����ʇ� �y���iX�h��^�v%��a���1U���܊���vb���jh��{g�.{Q�उAr�DǨ*[��Fw@6G<�y;�����Տn�![tEu�%�oV���&P?1Мٸ9��c�[K��s�U�����<�lP� _�^@bR?"IT��2b�H����]���%�c�
�K8���[朮�zy��Gw���c��`nE�`��K̒+X�T��m+I���ԥޅ���g,���Ц�HȂ����;�̣$��_�g7Zx-��N)-�U�yT���OW9i�����춨样�J�i����9~�)�'W-�V�Ļyy����x��Ю6�+�_�5��V[�C���U�I2���2���:�~� ��X�Z��=X��w��f��z� �ܔ ��%X͗UG:l�Vr���%�|���l,�i���*^��r���Z+���q���um)���6���B��2�����<ۣ��Q�9�Q���y�D����I�f�����k.܅&���`c�19C��}����Y[|z��6Zn�����"Cp�W�ܹ7�%�c��%�=�OU��N�i8'�������b����? �3�Ē�o�%��:����Dx��;�چ�<��{��D��8ԍǷ -h�f���w5�c�+��4�L�f�9,Q~wN� c�V�Z�ye)���B���ǯv�O�ҀL�̳&��^��%�a}�w[(1���F���3�a#���qX֟����(�5N��M� Z���q����D�xG$�p��o��Ũ�.����⌒aY7h�V-7vv�5���
ǽ�GO5��.����G�?DB�'���s��He��N����Ne��H��P�ZP����c#��,4��A	ʈ����Ե	�p�>]�Td��!��(繀���آpL�3�2�K�c�!(�W����@x�3`	ו{��<a��uj� ��