��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1=����V]?J�g�t;̀�<K�����}T?͉�F�([�$�f�0Ǝ,��,�2u5�z��d�����l��/[x?f�-&��� Cs����<i�KFzH������:v�F�[����?�&��q��b�Z�%�]�ӏ�@�NWǙ�="���hF`^xg��ϡ&�����C��o��P�>�dU�?��^}��5B���s���2i8�ab�x`>O�44D3bS����˩À��4]5�8���LJ^2h�"��(FO��J|��(�����ˈ`��T�'2#��ʯ?<J�fG��R�nf����S�Zc���M{��jfB?Ċs�`ʎ*ʶ��1dh�q�T�S�Xh�W��y[�11H0�mS8��I=%!7$P�Ǯ�� �,y%B�A9}V��\�?lSo�1uid�s�*L��{` XJ �7��f���s�3� Z��� 㖸H�/��<�lL�h
N��t"bTo��#i ���׌���C�?�F���?�_5���;w*��W��l8�q_�y����#$��`��|Z�T0�9�F�䓠���V�'��hC��]_������{�F�O���nU}4*QЕt�%�8�a��ݸ���^�4�h�Gt���x����6k�ށ�Hu���Ӹ�މ�#э�A��<�\��KK�u)c4��Z�c�}H�{n�W���2�T�i�ֆ{�W;mES��5lh�!�|��"��^��Q}���iya�e�p��So({ӈ��2dZ{�g�}�����~=ς'���8�-�@��0�g�	�Ik��Z ӁS|��9��bW�(4��z��So(��v<���O�f�$���6��]��[�-��"�pDA�1>F�h���֤�ŕ�Z\TWQ&o+8FK�4�,J��si�k���Sâ��ݱ7� �����;������Tc)��Tʿ�(|���������rslV�O���k��{�v
ɀ~@�����ޖ?��N&��&��@3�#v�X�[L~J>!1�Lo#�?S���O��Q�v'�
�$e�l�c��1J�%s��bJAIQ�A<�Z�?Q\�����E&���d�{2s��3���|�l�%6o;����x i����H��1�%��J*�eAM	M�=��̹I��x�� m1 y���wNp�����Iٮ���J"�tU8f	'��!ɕ��8��>]_aY�9¿��*`�u_s��q�Yt���%Ti{�bs�-���%�,j#!Ϥ�!��Τs5�
Y�����:�q��O5׌���k杇p��-?�5|��]�j^���h��./�rt�����<$���Ӯ��=���i�,z�X�5��tP�X���%>�?7ؕ�LUtꀼ�R���~ZE�g�z?V6RN?x爢�N���_��H=ۑZə%�m��WQM���(��h�b#U}�SY>��ɢ�����X���A�u�P�f����S���ѻ$�{_w���;o�������t�-�=.��mԓp�ʩ
z��RӴ ����mic1���ݳ�|��́USf�a�Q���$�Z��k��EtJ��O}��b�X-ze�y_���P>�uf���*ۭ&HЧX��������VV�.�G4~�ߡ��>�'Cr|E�!�:���Rs�߿���`��!������K��V��m��g8%�S�Q�q�d�ڈB�LI`d��~�Y襸FCa��)[��M����Cu�<-�>����B9^��w�E��6��`B���*�\�&q��~�P7��4��%�+���8sW�%,a9�FV���1�\&p���G���6u�Lw=�G�X�iie������?��P^�]�%�G�(�2{?�W/��Y$�m}��t��ÚtƘ�i̕��G���6w�Wx}�TY��7�bG�M+�P��Vi{��T��G|�o�z���;��P�$]Y����gώ,�=�X�#�!��v�
-�l���M���������V�uo�O�aY"�-��}u~h��k9��TN᪨�i�����!ʡ*�THF[��7D���6{�d��$���M�&&�f���h_L~�^�Q�f6o�籗{������Rͤ���I~�h�Zw� M(O���1΍D5��~w)	I�0n+�ho�XV�����n��`Wc��% �>5 g�@��t�QL�*}�L�<�z�IUi�I��~^�V5������ʍ'�J�/=�Uzhv�f�H��y�8��<]qF�u��h0���U'��D��ɀ Q^�q
C�C)\Ո���=4d)Aذ,Y�z���G4M���ò�����B �J'�Ͱ���C�!G�� C`� �*-ޯq�//��p��ʥ�x��E�-,�q��OJ�t$ޕ������'��'9>��M�R�h��悸�,��1K T��+8���4S~�ڎ�����<���љc}�m��kj+�� X�*��i�����ہ�����@���t�j#vF�0Q�@���/W�AW$*o�4�V��&KL?M�Ǯ;<j�����n"���B	�$��Y�t��-�@!����"^_����%��vR���"��m.,x���P���%��?m䧂��`�h�v�kh��d���i�o���(F�8��л�=���y���!�ś��Tm����������9?�����s��'$'?����y�|�5Pޒ��,0DC9c��1���u	΄��	��pĸ��pj����b�0�u�1*v$��f��;�a��MPZi��AlΆ�3m��{�R���,3�nq���zwk��|���̛M	���p�-~��_-�������h�nO��xKY%��b��@�ټ&8�Z����`�>�m�{*��̽<����-
��ҝ3�PC��'Ed�!�;7�����	�V6]������#h�wQ���.�G\���\��
��.O��*�9�D߀pM�V1�M�i�$Se������T�Z����l�C���FU�6f�:"��s��
�-��(�ʱ�=��M^ ]�@X� +	��'Z���׬dr��4��'�i�`c݁;)<n$�
sY�*='ݎܗΐ�'J�Uly����*BeC8���G�Ȇ�ٟ;l`�>5ֈ��t߾�"N��vu��-6>��q��wЕ��1���k�<��8a:�y�7\����I�W��$�)BĔz5�4��b�� 4��}��>���1���n�?�K��Ya�~!������+Zd���h�2�~�ETZ�����Wh㨬<N����f\�J�'�=t�d0bZ��l�{��=�
c$�ݙb	$E"%"Z竊������.����՘~B�q�5�C��j��s�y���Y�kԘ��D$���;�v���N�3N��q	<y+c3)���y�5�y���r�Q3A��";��H���>$O`�����0.ղȉb�W"~Aם��U�~��Zz�MFb�dl��a��]D�pq2�շ��t�h�?�w���'[�?�N���xhL�26�՛�Dė� w���ʷ���]\�q��a��h����c$��s�;Xwːuq$.�\�a��I3L��,��Y��<���yF����BUf��5{��!���]Z����=g�ר`S ���=:�T����<���SK�v�t>�Q�ٜQ��1�xsY^9/��#��x��b����,�;(�U��(םn�)�al��q��$������GYMO��pj�⠞F�ͭ�f@�ZF�V�5�i���hc�M�L����I�h�������ȕ��a׭��m��cܯ�)����6	N��x78��;�M4��RLg[�a�A՞�v$}���\�֢>O364a� ��y�R^��u�y �`l��g�3J3,1δ��}��m��ܚ�����$ߧ�J_�F�sM��r{�aT� ���!��p�p�gz����[P��QҼ�~&?,q�Ո_���M-� �^���Ԡ8T
��@�hnOɹt�@">}Jfb�N�+.�'IV����9�������W�-A�b��Ml��7 ԍp���1?�GC� "�(M5#-�8�5=5����B�UpU8�Qn�"��t!�t����8l;PO�9�`�u�|�y�}V���y�e�`jFu��8~���,F�268M��6�F�"�aX���n\�ab���I�-���y��eB��X�Q"ۚ6Kt�dG���ʡ��~���4���H9R��HXP�"�,w�����;��E��\ ��h�
��o������9��iz^L�oh�n�p��Z]��`uOgtgs�o)����|�؜ɅB9C�@��l�T�I�&�U�hf�~v�]Z��{�̒-�lfv-���%�p��f$]jP�$1�Y.�!���ű!��<��%����n�d���Gj�4��r��]C�A@u�40��W��]�4+	`ykx��y��ڙ�ۖ֊�p�#d|% V�j��S��E��ˌ�dW���9��oW�T��(u~��{�y:�m%l�8B�m�GNS����&��	S�쬴J�o�����{�Oa��Mv�Fٵ�9���%ީ����6�蝣Ūk@~s���FN.N6c�:�6p���o�3=�C1��ŏ��T�W��H�⃟�婾���/�Gh��6���+F���ѷ������	8���9���aqTz�>�k� ��ܼ��m;vɬ���H��Z�ө/��
�d�`x3�:�)7�Ds�� �a�>����*�P�k��W���_�n��8�VF����Lg�k�8��~�w�v�@�A!�1�H4)����m���e���vy���e�w����Xu�쟡���g�:���Yj�|�g�"�8�Ij֌u�~,|�M��]G;�ݘ)>�b��C����
���8�i��� ��ǖ��U��Ek��.[Wr5��	i{w�\�qh���x�I�V,8�A���e��#ۧG�ew+f7Ȥ��T������C��jH4�`�4�6EM�
��V�����/RPN�t>_�01�	2ű���Ш�
>)܈�����[�:�����$��3#u�e4���qX�?���l����1�<�u*��'� dztH�;nsJg�:)���gڼ�$�D��b� �Sl7r�A�.���Ӵ��a@�����*��/të��ۡ���2�7K���,��־p�\#e�#N�'��~(4%cϺ�#�W��鿓��rQ�c%�B�h�,Õ�v.�Z��1_�������Q�Eۖ����@�a�p�2Q��\�EpL�^�*<��Ԏ����{��n���Ƽ=���5����B��-��t��o��`E��|����T]~P�����u:Y�ҼR������y؋��g�
�h	�`���7�]���"J�[\ύ��ހ�"�^&�#^��5�T�6�V�¥<�)(?�@;�U�[�!����G��C�s��s��\X�\�&�4�S��]l��6�J����-{�~8i�*�8+�NvM�	�K,!]ݦ8�����5A�{B�ls��ET)EK�p�X
Eq�-��X'E!�jjMh�|͊b]����qM�sS���㯱I�q�ܮ6p�&�F��Xܜ�F|^��$�ʏ���%$(.Rz��d�4��)����Òj���QYZ#�CvdH7�~��YX|�ՙC�uCD[���]��~,���N�P�흌G�2= D�?���l�D�����#�4�������n<���z����}(O��*�r��ճ 5Heb��p��Ujh�*�����yO�L���ط���&fx
�Uz�?��l9������W�������ޒ�����'��-��ry^?�F�0S {���O�=
8.�ؖ�~'�ލ��+�O��$��?r�0:��8I��n�W��n)֋�@�$���f���a����g��s
��E�B3!��_}-m�|����
֍��-�
SjuZ�k�@@z�QR�2SEQp�gS�260�ۀ���5h��Ur���X�jc7�6���!�|��$���v��*&�W]�PL��0�� � A�//��J�a�-��v��5�}�I��p~�B����%h0NC�p�GdrX�����V�����b��q~-�6��c=��X�U�z?���Ρ]�#v��=����,��g��v[�=�ijY��|`I;7!�F����Wj���Dd��K����=a����q,�-0�B2o^� �7\jYEzb��>���+��갓?��������ʺ�Í�N�l�6h�RFrb�a�9)DG����#�F=��1��.~��!��~���s��
c�lk�ޙw;�rZ9���_w46$�us*�V���g�C��S�N�"��ru�ѓ`�A�Z�3o�ň�/Y�<�4���*M#buNi6b�ޱ2���V�4�\���hlO8B�n�E)�;����