��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ�����DŚp`��G�����D�����}��s@���L�D#�� 1�O���:��ԭ��(S�K�����qG�k�: �g����A��k^���%�0k
%�����<|�m�у��+�Vv�%�B�%����5�n�vf������'nZ�Drd��C��uR��%�`��"#�"HO�y�Pq���~Q ��C�5�bN��w�y�=�v䏦 ���M��䂞�]+��징�����!�yo2�,f.��|o��e9��F�����4��<ٝ���R���P�
snU NA�-F=@�C�zV< E���F���?�2��M��$�鱤��Pj_{�Tĵ�۸��g�h�]0����"dd{PT��d�&���fb��;B�d�i-F\ z�6�q���)i6�h��*��9�ln��n�O�pVޭxN�j(�o�'��4_�����R�Q���m é�:�z�M�\F���4��w�K+����҉%�^z���6#	��J�u��!�y���c�����}ȿ8+3�R�9-���~��]�`�=5��%_�f��Vf���w���0$ �,�\�52aX�	�D��/�����Ш������{�j�^p?�^��oF�l�G���"<�AޗsQ��Y��2z���c�M5�0�����@+��A��4��
�8�����v�b"��l�����4��rϻ8��;�]L�K����X�����&��.$qy�S;�	Z>�n��}Z_�X��(}�<���!���оN��:^�}��7
�-v"g��x�jk0��!t��ծj�Ӫl3F�ح{@��"0ݑi�l~'��4�FKe@�_� H��h��Z���-��0�f������@�ɳ�(�־b���*������r�@�n�]k�HĻh�>EGL�x~tp��?�>~�XC���m�hv+�خf7 Ro~�s�6������ 5���!G[��F��+�L#i+������+,��F&�IG�P��+.a�Yd磒���ޠ���uD��g�RY9y���8�cS!�kl��m�a"�������2�N�-ڸ�r���<�]�yf[RZ�s F�B�f�		��`�^������$dM~�{��=��R9�|�T��cr��
��鉤*Pd���"�ʀ8*w����X�>���jgTg��'Ѷ�ώ�:v>"b������o�1s5g�+�M�%������l�)(���
�g���l�-����k��YwA�Qz
�Y�6T������熐���i�)��꿈y!���ܱ�eN���F�M.1�Z�E�{�v�2p�=\�W�~A�DF�4��뫇�\�r�n0�p�&��"	��^Y�b�_)���ػ6<q��-m[&R/��q�j_�Ȑ.���[P61�NߓhB�������rA<^��;��p�6uǵ���/�H�	��筎�W�_Ȧp�}$.#�?���R�(��o͈e*�kIM#�>J��s�ڻ#:~l����V�µ��אΒ�����ye�e��{�\�ˇ�R0Y��Y���2�#���H�����'�vN��������Iz �2QXʥ��$�Ai��V�K~o8�>��J���)��*�o�.����󣻎9g�)��0�ņ�;8S[5��meLԷ�$��Ƿs��Hp�2F�_������5R�=���~i='W�ks瀫'?Pظ���}��ɡ�v���,cl9"P�t��io��*&��Ύf�J�aK_s3��2�Y0j�Ix�'�YiY�ZǓLLdPo����W�H����ځ8Q�ⱌC�.��㭟�7a�#�w�%B}����v)r�J2��c��]=Pԝg9;�p`	����IY1N��$�������ּ���z�vz)Ω�c�ٙaҸ&����
�Bk���<W�d���ipB-m�脞|���'��>��'^���aݻ�H�5����U	�%��Jmj)IE��к���9f��L�ɻt�@w|���2קM^��	l���/B����e�}K0�;�]�� D��c$���b��X_���|��=�x�}q��;�m?�� @M(w��z�ڋ����Q�b���,{�,�a0�f�M�H'?�G��3��8Fc���]gP��x��`L�W��IR0������-�շ׻P�p�y�.���S��[`�C���Ɵ"�	~G�%��x�f*4I���� E�k�*\�|����WR�����:�ü$w���kq�s�{@,�T���L��dM<�t��e��;�
�����5I��)��G1'�DN8քª�u�;8B@�B��-���`��-:p+ca�u3d"m��䪯k�R�>A�"�ArLJ߄�&��|���T(��L����x����
�f)L�E�'�����v��<3�A��ﻜ�`���q����ȩ�H)����G��(=t�/w�$rҒ���ˉ➅�$���[Pw�h�b�}������:co��h��|5д9���4�7��x��[v�(j��k���k�I�)�2��ך8��(���#	�C��\��Z �Os�i�Xl���m��qR��5�cװ=�Q����D�]nȷ(Ic�]��
���n.ʹϢ�43yN)�1��ħu����}�R߮ۋn�ʋù.6�MN��8��w;��P�C���M~��,� Ʉ>�ka�Q����z�����Y&�#,���$`.d[��Jj G�l��HN�l�7cd�S��	m�gr�۸0�J�+��/�HW `�U�s#�H�'�,�'3�x�(D�q��|�JJ�!D� �t:���f��N�eCXlq�D�M_������!�N$��Q��b]!VΛ[����x7O)�d���j�d,'{6�l^[DG�����j� k�m�r��?�5������c�T�J�������*���V�Á���[��I�l��46D������Y�+�E�\���rd8m��#�˒G���L��[�sD��k|�}��[&�f��b�ѯ�WV�e���*E�5L���LXO��6���,Ps�����`!�\�h��>���q�
M4�6E>�'��㵒a/0�;�jٸ�~0Ih^�j�G�^�jy��K!�ϬvBrfv7���S5�����I&
�'T���[��f��I e<T���G�g7%1�/�S��s$T1�A��X�#�*��e�P^��\4yFe�[��<�/鐣i]�Ql%{�l����;۫�f�.[z�sH[��A�V�?��ي�M������4pK�@�e*�4nBG�C�n����k+y>[Q��9b'V.�
�H��"é���@b��R�:�|Q����+�1'\�?^͒gz��]�!�̯��\�gS��k�:��d.31v�z����+͸��VȊC+�u,�]��ځ��H�5����c+���A�bդitD�8�U���3���7��^;i���sIri+`g"�rN|�Z����H]w�ݲ�z֍�H��F�E����!S�����<&m��zZ�a�0�hĸ�osM��F��R}dD��*}�5/$T��m��k�IbV����4�3��ؿ����inن-�N�֜�$��I"�-*�P��s� k���)&�d&�R�_'�VǺe��k�ڔK��2��VǊgB��s��䂙mDVy���y�P:~�"a��=-0=���?��2b�{ǡ��zb�a�Mw$��Y&+,�[�A��X��U��5�Ζ}}ۄ�+�D���{wQ���5��oׅ��D1������إM^�W��qƯu~���������Q}�'��<��O|tרI�n�6�)��z(�!����CU�oqTX�jx�9_�� t����:&����\��$-���Byk�L����~z/+?�%��U�:�E/��mr�m��@�頯�EUUπ/{����V@B_�u;�_��R#q�(�'Ք�"�G�Wb��|�(��Օ�噃�`�+&Bp��=|q���	������ˤ�uG7i`��Ax��������j'�^����&0�C�m�;��N Fk���k��/)	+2b�M�(�����O̹a�����j��5$gH<�nn�W^q��sm����H66�M�*�����]�\��ɋsu�0��� o.�tesE�^v}���)&���m�
ϣ��e{]�AV�n>5�6b�Y8-߀u�wp�B#��U�F��Wu*�~7a���#&��Ł!\.2	�Ҿ�����R�	�~T�-M�Q�9��I��`N��B�2�+��W�[fe>���^1�͎��~PەA�~8O�~6'��ҥS�G�;,�(\���6����s=k`�����.��&���� ްXr
�M?�_Y�jy�U�f���R }��h��I�3��@JGW� g�'8�$owt�Q�]�yg$�P��>�z��q,�\v4Հ�pXyʹ�2U���&p�τ��Be���Ms���d����H�8U��h�v�R���̞Kl@DKz��m/Ґ>�#�c�^ᦟ8��iN�.z�4ʗh�ZԱ!T�L�A��!����p�����Ŧ5�b�'�4�Df-!��D�\wAԹ�Q���Nq,m�B��������+֬�����O��l1�p
ه��R�-`�NgA���c���'��TuJ�ȉ�O�ƿ��Ws�M��Z>���u��3�yTƌ)Y���5}-�mRgD��F����j��2MN��2���)���9Uj{�9�0����R`�K$�	/�b�����	�$�Υ�������c(�9�UP��%��^�A࿍��ɛA�fj�j�\�Ӱ�f��s�y��6Ֆ����H�����x �G�^���\x�q��L�'aPG]�����\X�E�_j����,e6
q�"w$�6�k��Wj��z�.�����bi�z~���y��$~���c��%��o�B;�`ΤQ�����)�4$���5�bi�er�a鲫�o�}�>��5���yR�t������q18� ��Ȣ�c5=��\'v���ɝnM�\��Z�[�4�Pi�A�[9P�ks��S��G=g�w���V����H��w�M�@Ǝr3]��6�\�Pp�:.�(y�Fs���1�C���H��Z�fѱ��&(���be��� �Uq�.�-!�nVa�@*A���Y�{��MK:� ��Ln��[��f&S��:�6�Σr�V�ۇ�#��8�2�BG��������$�"���~q���,[~8��Սc�d*�iυz��u�Ɏ)�5L��������+T����}�_�n�Q�9�Ӂ
�� ���;m�O�;R�EPP�h�j"F�y�*����>)hv����͵^BKEQ �)\�O���'��!��e��ڧ��SgL����-$eѝB��7��ٵ��E�*e��,E��a$u )idM��v��)�H1�\�<��Vkhʄ~�
���8%�K>l�?6��b�^%�u�_���r�a���W�WuW���yVd�j`�,����I	9�`��p��A�;XX��	��q�T��Hɵ�m;�)�<v@�|����m�#�<�X�]�1l2�K�:���k�P*�\���\�u?����v�)^! �x��p~ �BEƧ�+���#�g���͹h�B��[Gj�VUeA�f����B}�A�M뽯�%V|�㜞�'�e�E�t��w����y����f@�4�>CE$����y��*4}��W>J��!!Rݫ�Oi��x%3T���MT�!)?���<S�"��(���k9%�\q.q�;��ŏe<0��[��2.w�A*
��J�U�6�j/uCr�b.��L
Xw'ѣ|�CkN�JH3��H�P-S:&#���|Bj��� A�t�IR�j(*�hX��T{��RڎX� �Z��r�)!���q����q�QSaP��*�0��>���BYj]��4�_2�" c���P�5��l�;��#2�&10��V�⎲���_��;�K���Q,��d=���X�߇U�h�l�3=��}ܔ�K��4)L�%����O!o��(�3��04����B�)5�<�֍ظU�U$��ʃC�>��ëz[�--F�Ϳx�^eRER�v�_��"{|�G^��C������ع�
��x��%�h#,�-�8���t�S~VB�Sus�V�t���G3)�M���F�������B���厏����)J�C���sg!p����~"/K����Ԑ\kxd\�oDZ*��ZwՈ�
��9&��{bH�x��L��H�Ç�����r�q3i��47��F�u��~n��\��q���������w����ujH��(�GĠ�g�G<�b.��<Q��|�X騝YA�J��Շ)_0L;,���@�t#���l�fv�,Ƽ]��gTя�m������B
o�Ir~zwT=��U�9~�Ę��}��ų(~u�����D+(���������ݱZ�WRR��]���E�:P��@�SR:��L��+/�
�H���c�(P_�O�$,)�/&�K���vS��c�y_	��n�L�:J���=S�Ѐ��S���Z����`��&n���n4�^r����++3�,>el�:�D��O��4�ё�^�u��Hu���(�K��i§y1�n}t1ӼF_�����M��f{$�C�ۧV([&'H`Q&0�%�~����Z��么�k�/4�{��_����v8�9�J��uz4��y��=��'&��7�UU*��ٲ���{}���LQ�@Ss�Tu9fr�w>X+�??����\�N�S<��O��c�q�SY��z3-D�g�R�doiZ�PG��"q�p.W�Z������q���ϭ�JR���9QJ��x�f��Nh2���
�.(���Y)#����{�8���U��P��֗�n�8:��`�eO.4�5'2���+x���1�C�4�s���nA{��#�xB8�ǵ�V!��)��S�!x�)(���/��^N�mG��xp�U[�|^�o�+H��io�}Iv��;����R�=�9.�7h#
�7��� ��	��SLi���R��������\��q�����z���)�FJw�m�0bw���_�U-��ec�0��v��K1�/=��7C��H?���>C�!~��3�=�Z�6IB�s�R�%���Cd����?Ki)F���������,�}1��X»���tski���A�H�L��SΒ`m8b��â�����5inD8SvbYƱUZٝ �����_�/	����T>y������^CϨ/jՂӕ�r�c�&E�9
�}��>yVC?��,�=����>���Ce��E��Ú�$S��ڞR}����.2C~��1z�]�ɟ^��`�Xy�^6��fNg	�_�R �q��.�������<� o-\z�޿(n1�w��Kg h��)ܴ	q ����dW��7�*Ѫ��n��4�B�D�5V'����ir�Z}V�yu'�O9���󖎸E�Y��`3�-�&���b�=��͇�ّ�~�¯�0�"7m|�XT��A��b��
Q�.�ٍ7)/�O1��,�{.�A=��4x�lda�=�
A�OHkӊR��r���D�I�\��v��V�a'N>�xc
�.7Z�����#z *U��z*�����`a�?ş�1|�=�J�HF��yB�����zf���p�Xu	;
�x5<���k��AK�hݨ�,��d������3�Z,Hs��A� c������oy�'bc2��I���.H�0��e|iõ��f�nX���ng�[���+�ԹY�]�԰_U��+j��bj�>�eJ{�&Bo���6���,��.G�k_�%�x�����˽�/6�Ӿ$[��^�kqT�����Q��r�ݳ��OU��x��=�L�2�p��	ɜ�p V�X-E�Q}u���A+��`4Ou Hʭe�PF��1�z*�U���-�����,�ع�W�6g���U��7�ZA�Z�n����Kk�mǲ+����C��v�v��	5O�8��;H0Ά��Pbl�@�d�Ȝ�6����򃽕��\�B��#�y�+��߈��c`�oi¢f�b�X�q�+VF��l�|���%��19��N�%����b���n;�D
�O�&B���g��O���`^���P%���]�(%I��2KMr:r�����&�!�c���n���b�68�D*:�.�Z!�`���/N���J�/֒�H��r*�:$�)s��) ������*�KSG`����jЦ?$;��1���t��֛���*\Ȏ u�egX*����9hbF�1��󽬷�t<pj3��E��>�E�_^Y�w�.�������_Gj4W�W@Z��Y@����O�r=�B <7��m������(ى2�g��f���D��
������9�,���$��ca /9BZUi]KH�p>��f��"���ݲ3�WhH؜qm)'���ǹ��R��ݓ�z��gΙ�C����t�M�袢$����=;�G�����^��rJ7����r��q�t} ����wbe�� v+W?Y$�\�|O�ή���JHڎ�m*k��8T�tz9!�y�V��}\3�;F٠�F���hl�냺�U�:;`��@������Ur"�4���躹���;���Z��34j������9fK�z���~�a��b�o�)��O�B���0�e%	lc�3�K���Y]T�+RB�W@J\��a1��5L�bˆ7^����l��1�v\���*�sH�0�*�1T��'�U��_�?so�a��"�􎾒��D�m��T��wq�j!1�C�8�A2�����X���B�[V3{5%b�������s�t$+�P�Y�W��/YfT�L6�*z���_�I��s�M��8Z���P(٘��]�>FΕOO�����|�j�5M
�&�[���k'�c�F��K�/��8����"ʺg� A2g����T�doT5s=l4;<�4ߠT���T&}m��Wd���V�knL��k��7GF��Z������рJ�\�F�C�l`�R��j,=�T�>;}��1�L�!��� ����O<:�����-O�O
�h3�H5hm�]���
�D�<��Hl �����	F�J��z:�[���	�0#�h�(��,�s����Ռ�F�D��� ��eJ��.>�'��g[+eDF<��O`[�3iP�
��[@"��b�� ����%�M�n�🫩�����f�jnTf�,.�?,M0�t��D`
�Zx\�97��ތ��SFtՙ�\é�v$��?���1��� )�H�O����W��Y�X�މ�䅼��yb}��b�BF!���-�v.����Q	���F����Sp#"�)�Ý.P?0\?k���s�!;���Ia�zٿ�5J
�[A/����d�����謓����@��y��Hn�I�!����2�� ��1�J[����G�˰q
^� c�ѷ�J���.�'��R+��oBӶ���} �.��c}�m�\�%H�M}%Gx0*{ƙ$�1��6J�p���0���ۚhr%�e ��0ˁ��x2K<��ؒ�h�0ȑ����뒇������?���&V�7#��ʮ1B�Sմ@=S虅�{C���3w6(}Ʉ�!ł"�Z��73'�_�}�*x��9#��w�S�VX$
{�����ܥW�D��p��p��K��-�����*�Wq�.CA�ȉ���d'�q�ChEg�"�l��(��~6y�������̃h�$B�.�S��7��N��^S���ۙ�,�q�ê`���jҀ�킽�o\���&˰��/�&���~<�l�SWlc���ū�rŝv�T���NN��
8��t�\>5A�D�U(ٔr8��c��wr>U���ʥ^���R^V����s��u�S�� ���^����%:�4$,�*�׮P�l�RP~��4���˴��Ro� &$�O5�?h3��*�d�Ƣ��ʴ��?b��!�a�r���&5
��:8�?Дhֽ�SH����u�kOfeH���w�ί�a+)L�؅m${�/_IK��;�()���9��z��Z!�,� �:�h�R0=�	B����ZO�)�O�E�ݞ���	��r?sըOA�_�FU�v�Avg���M8��Q�e��,�P���Oi����O�*`�H�/�b���}�(%]�����DRǇ�c(��,��TK�,��ّ���ɴZk��h7���fxR�B�S!M	Z��F�[����s)���*Iy��z�ze��k�p7##���,��T�qx��#}͚�}��CvU�Ċh������L����s�w���@Ny2O/�^
�2T�WXx���ǩ�������"��A4W��Cĺj�~B�D�1�B+I��AYmN�j��9�WPV-����������l<�Fa��>9v߷�0�H����U�{�. `�<JZ*��V����ӂG�:f���Dp��P�n4�>.@}m
m]�O*��0 ��ܻ�Td���V���1S5v��K7j
��w�MӲ��wB��V���O@�b����h0W=�&�ԣ��'��s?+�D�5����&�x���<ɎH��X�4ۣ��$HDd�P�\��r����@#���ב9J�r��,��C*鼃y_�i���:4��i;���u*���9��(�;�����Y+4�����KBqHI�Z�-Mi�=Z��k�Rr�߼��</0�>���3E��D%�H�%p�G3�7�S72�=4)��wmv/GZA1�S�HZ��Rv�ĭ�H�6ry�O4Vc�h3@�a/�v΢���	K]z�]u��	x�����(�%c�jl��_n��e��̀��M^��0#��'��-�ZLU�N�<��m��?ɰ���\�|�Ƃ��_}zg�����E��饺���lH�R��:IJ�w���}%-`��yM��%T)����,��"�Г����QR��R�K�i��(�ez?_�|=�܀��F��}���*�Ph������qŹ�+%�x��pn�թ8A>;��ǀ1�w�m��p{�f��pKB���,�r�Ĭ�FP��I����Ւ<�r�>�Ot�L��;�*:��]�xW;eb�g��M��N �ֶ)�D�kå���K�ܓ��˿��qW
Z
�La�FvD����f����0�MJ�\J�_��.!����r�ص�X	,:-�4��?�6�ub�3�y�z$;޳��Z"�m,b�5�7}Gi�rG_�i���R���I����*=�g{\ G�t h��"iwm{O;��?`*����~�S	\Э���+�EI�ݎ+c���Ɇ8S�T�^a�>�٦e�aƃmV��Zk%1Hg�9��Q쳸P�.�`P�@��T����bQߊ�4?hС݂�A�vE��Ex�J`�g�s���e��5I�;�g��lu#���q�RҽH��p�