��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ�E3�N�j].�uj�A\3�/ꤵ��W-���߾d屍#Jpƅ<ysR Y 2x���lFeN��q���R�����W�$l�g�kL�ʘI�ᗨ�ת�<G�7o���3p�d�T�8�,�c��dn@7�����	~�
5��uc3��9���_�#�z��&�p��g�Y���'�!|Uh�O"�uK�����}WU�BW�fPh������Dς��Isx&u��P?��&Byi ����*�cPm3��\A��}�l� �{���9,�r@*6�QDjJs��%^|p[�H�lٽ[���&�i�,P����shr��4~�PQ�x�-&M�>��nް��븤��)@$�x����i�t�̤�i!�وޔ��2�/� &�ս��+x�͍"[���恒���jw���%֏��I<"���m8�cjg��Ϡdͪ;��t����<A�"�?��󞐒Nq�����T�&�t�Aϓ����11��ՙmn���S6����W��8brჵ�_�RCڪŉ�<�cP`�w�I��PVy߬����B2A?eg���n�
{����<��r����$&�ס^y�g�_�p�ZC7Y�����)	n}�|1 �b&Jƌ׊��.����GO@�y�'�0�~�G6ER��<���{&M�'Л+�U��ӭ��W��1u�[�kcy�MkՆ��;�4��	���Z�.Z�>-��7���t���K͆���{y�|��ĝE��
����(��^��7i�f��>Jb�h����˖:�Y(�i��x(����0�e����5�"xL�ƹ����8��O����z5k��9�{]�1�������	:���B���x24K��75����;���x��K��5
�8�k�X̩J��]�}3WK�ú�$t}O�P@@���&���,��/���J/�{i�~�]a*2&�hyV����h��%�hC�̓��&�%8�fX����\�;"g�[�eq#��i���-}�
$ܐ�<�z)(A�nwv�ހ�z�����'_Dc�f_��?�&��6��s���N�l�F� �.%X�k3Dն�z�vc��X�F��lⱚq�V_#]�e%�(oH�+�D`C����-yZ���7��������K~=tp#�@"
I�B���;��cB������WK��/aoz�?혐�!��n�@[�
�!o2^Zy'�@Ɏd�I��`fI�転����Sᷗ|���EE����� 5S'�7�h���Xj�8U��~D�c�`�>��<n�$D�7���#� ���H{ixe|��ХT۠��.Ҵ=o)�
�Z�*�1�M�x�a�=p���Q��^��Ȃ�%�d��Hj�1nX�=w�)Y*�T�Z�w�z���C��2Bj*Ъ�&),82�� C�o�����jX��M	8�Z�nZ��z.[���\�Mj�U�� ��%'�\�J8e�'f�-H���v��V���X�"E������뗓.�;�S�W��#x������δF�7\�Z҆>��������+����jJ��|}ہ�P�#�� D9D|T����H�Q�>�.wg	�gt��C?�^kP��i�����0���D���ds�"�N)GS_5�y@+%l-2+��������R����ɀ�D`�����!{��#
�8�FT�8�-`���t�)�2�k��֒�Q���*-~z�6�gN���L�U�	�9�q7��~��P�ǩ]:�"�w�4��K����%ֲϿH��8��,e��������p��c�s�N�y�c㙑��}�rN�=bN�Bݬ��ۨ �R=�*6����Uo/=}�'�-�<���8rSbNN��S�'�6�r.����L�-���I*��M���l�zNi�k�
�e��@�5���@3���e�Jf�D�!��W3�fەU�ɴ��a���C���0('��&P�o|�����L��^n9��̕]���3�~���ԡ@al���Z�D�)o�'�nMlr�䛯�f��؈lr"I�B�̽�,w��%%���Ib�Sm)E���T������7
)GBڂp�-���-e9���M��H([��9���_���k�H��-v>�y����@��_���-0F��
ٙF{�-^���di,#���r���"�+�@t|ћHha�^��I�0��U���Ա��D��E��'����M h;��p�=
�	�s���2��T��P�P���֧s^I��yq���J����ڢ����vW%k?����ކ������B'{ᘇ\�����`$!R�I�Ek���t�YPr1��e��ݏP�$�C2ߍԂ�X��c���� �Y�Vҡ�njHy*mOX�*m8�P�����䈵���_������`��J�	��C�o�u
��a��n��C��i�/���OsK�82�0�W�'��f�<;������0!�D�	p��G)̔������.���E�)�=cm����37�z�F��)��k�P��W sr��~�W2�~8�����R�;2%�x����� `�s�ߚ�|��6@�26WH��߰��PA6���z���6%�澟#p�X0�`���`���X$O�� ��i%�&�+������!Cs�Q��9�68�Z(ځ�7�Q�4}5S���J�@ �!Yi����-O���kEU_��&�ET��#�W����y\~%��G.%�YT�*N��,r�Lg�R�O+@Vs֭w� +o��d=6�_S�m���8�b EF�Ϩ$|�ىִa��Բ@�Y�U"6��<���F�Ãd��5/�3�_�!l��x8+#N��pޮ	��0�X����V��Q���ۇm~,g)�� �g(��5<���.Y���#�T�f��n)��_'#D^<@�����%�U���iH��-Ŏ�$[׷����QI�g��ȵ�<\-�S�_CY۸(
�����x�v��]���a�����
�݇6梦(ݍ=��=�YC�!��3Eָ�ɇ���;�T\eekT�	���z�]bG���p=���<�ެ���;�|������ �9�3RT�aK�uo8i	��8��4������ b��3v��7��ն���aK�sw�#�b> /̥*qd�^`c	�\�E9����C ����WȘ5��4O������")<B���=��4|�[A��^;�"M�J�F�����x��m;��z��6�)Z5����b
ڭzBh�y�c��ENDB��KK�ǒoF>5�t�g��V1��l1���r�(�%�Q�H�m�����"Q�nK��B7�~m�Qʤ{���>8���oF�x^�2���(��p��Z}�a.�>��G��wڻ(`&��M����
N��_��F�g��EAr	���C���?3a[A ����^�g|�IHN=�RC6��%)�R+2$L;�����銘�j��B��G�1 �ß�2��{vdr#`a:�R���h8e��Hu��%j�+�A:ʁ��Qjx(���p�G�>R�� ��^6�J��~��N�P�:�KJŮ�~^@j1��5��ݺG��̧� g�l�y�x�)W/U+_���!�fӱYP��r��'�3/��ٻ�1A_M}Y���Ie��4����%0d��)�'̊ �R�X>w�V�1�jI��&횾�]X���F�� ����K��L,���V����s�ح��FJ�W���0��Q�c�v�`5��D4R.a@��]t��0���>S4�Q}��AYl�Λ(ܛy1v�k=k�5�B��ٚL�f�9sfƽ�ͣ��:�u!"��Y�����<az��3��S�(_կ$"��`��w6���ar��;�"�7�W�L$f��kb'�|c%�m��0��\�@֖3F�T��*^���\���9�Qq�y|���I�IY6��[�er�KB�����7o\h���q���k/�&�I`�w�F�;�=����1����5�j�
H��6�D��,�үPo�iEl2��	
��@�3����o��8ny]P���3����)2/ %J���R��؝\�_"t,I���Y_/iy9�>0z�`���/��'}=|{�Lw� �MSӪ�1wl���d���E����*)}��9��?���~�EÄL���t�A�OSd�"(�UXN�q�Ζ�� ~�3`g4Ew�>�}T��.+���
5�X�;��
2�����)�:Q�K�[oWaf?�uG��dQM-������{w	���:L�f�;=�zՙ1%�J(��Kh4� (U������p5��ˤ�(u���[���p�*�%����c�f#ĠA_���O�}����eP��6��7�ʸ���������aS����������K���)��"�όch�#�^YH�i�����P�r!�հy}�&�o�!W�
�ȡ��jtx�z$�@ B�F���}|G5|����� �R-���>g���Ŗ$�'M)��`��m��m>�<��+l( F%�j���J���NP��4����<{l|��G���v���櫞 W��=���l�vϝ��b;4Sb^�cH[��s��Z�ԟ�a$��+�tb \%�5/0c�7�\o8�{t��3�W�2^��
[�^�=�ѱ�F���}FeEb�m���&��8}��������3Ԛ� �r�Dڻ(k��Zg�S�������Y��DܱV�ng�h�T�3��X�솿vd�=�Ew��=	Ճ�{�_v�>�d3����I�}���kd\o��.�La��y3*��~���`ei��Ь������LY���Y�u�� ��Z���uIՃ�@ƴ�U�XhFZ��������z@M͗�1�8FН����Q�Z�8���p	��X����n��D�o���^_��4ki���~�l��x�DKl��s�?+2<bk7�ӌ�����"ig�H�x%B?m��9IO���AU�J�E�)�?̕~��M��Y	�%m	4��,,VI�	�Kn0B�8&"����;T>\k��߄?K���8y+VO��d��y��Z@*�0���?�o	\<ʕ�R�w��.����e5����b�
��)�ͩ�! ���1�3��m��*��I���7äd
j*.�u,T�p>���5\n�F�7T��c�W�7�É�)��"1�+��y�G��!���b�����rgW5�?K�5bP*&��W��㳧U3/�.��dR���O�����acF�B��1vH�R�+��H61�T�SLj2*K�k,04n� �x#���
�"����8�휁bt�զ�c!�ǒ _I�y:��LC�dau���d��SC81:-��dR/)Z�"�E��%f�@�;���,ȓ_/��)��JpC"1R��!)b�4��̿B�����;>t��o~�~!㜻~^v����)���9�0%����	�j]\��-kz���d/�`��>�� O�����Pk���r�Ep	�@���4Nn�w��3Z�h��o'1�GF���d�~*�@B!,��䭀���Hh�o4�1ы���m��l	VK+�b~=}�r��ev
w�Ǡ6n�g�O߃88�]��훸��l�����}�g����;0��S}+I�G�+���M��XG �d?��ӆ�)壗M�=�>[\���06&յ��3ș�ӑU��F�����O�tV\�*�.��8�\��s����P׵��Ѫ�����)v�Rf�缃�@�Z��Z{]�lM5�/���ajgN��8{���omoD��,Wр�ѯXV�C�o���a�4��l��N��=��'`��¨6Vp�+��4�]�� C�j:V��ן���_��L�o)db�x@�̥Ն��1=Se�]@.,!Az3��?�ji��3C`[,:1#1�%���z�	E%��@/R /�d���=�T��#({������Y�O�}�c��fh��X F�����g�Ws����r:IJ�Q�(bH{�O'��<Aͭ��1������{���k|~L zm��, o�.�M�.��8��B�D�RFN�'�ՕU:�> ��C�?�K
���ۦ���YaK!Ej�&N���it$��h��Ԗ9�>�bp�u5_�����_>*�wy|��%��!���h��� y���q1��7��X����7���~j��f�9ݜ2D��g����.#9Qǆ��P|,�F��j�y$[7���|���d:��ʘǘ�3��ZrZ��@�_�]��J��Q7OK��Uܠvӭ����>�-�=�z=�Ͻ�`������	�c_{�ة>�`>�^��Ua�à1Pb�]O��a�B�` ̷�c����F��W+a���E&���BU�G��¶�,&�JX������#��Bi�.q�]r���}C�9�E�2�>�y<*���"����4�BDp٭�4-]hްT���x��4�52�r����'���C��=�g���>]�o&&�^��?*l���E�Ke�/�BP��!��^�wia��[f�\ {����a���+&�8��<�~�:�ʦ�]���r�[�)Nh=ч%�g�[I�����(.�4�&��Ƣ����-�ʤIڭ#����[t�΂%$?�X7�e�vMmQ���X#B�e8M���"�Ї�m�\�CL��\�p�����V�P�)sߏ���������δ��z�x�b� Trs����;D���'8vMHN��b�.�%/�Q\9�kG����08OUh0�VϳP�h��d�Y`7C��3Zv5�ܮRǊ|͈�mP'�	Y��f�X��.�M��xNK�Q% %��<�*���0@��������=�a����<N�'�B&�Ϳ����cG ��.���`�+�������Os@�����V�>;���U<���	�!�S٧�~2 ����WS��zy~y(`�j�[�;xW�>���K����0��Jb��u
8b gᏆ��I:� �g+�j-~�kD59��r�,�.��Y��WSS,ץ3���'R2�ҍ+���,���T��6�f���̊�l����I�C���i�t.؛�a�sۥ;�������=�N�ɓ{9 �0:��kIy�{��_"�}���)�E�����H+H�Ƒ��v2!ʳ�`�S���!��3S`�f�gOy�x�0u6/��Hr��A�&��&��?@�@G��B"FB$M���.C�S��Ht ��$�9�6M���/0d�	�'��ך]�Ec��` �c�`�0���U��{���o�&�.�q�e��{�T/�:��	Tn����� �Ym�6#?˲١�"r�����Dv?�d�9���I���������Z@�-}�3Q�ħ�{�&mc�Ǹ�t�q&�1:�E�9�ťO� ��A���ԧק�����9PE��f4�h1�Cz}�7� X��X޲ ���t����9�a
�����XhگĎ�x�Q�������[;�����f�q�"����V%�JvA��Qd֤��m��$�P���gk]9|G(��`*F�)ʑ�s�9��ݥ!#CI仧]�� �`��ey?3=��"����bN�h�\�ׇ�(#�?���;W�X�io��C�Y���L�5Ŀ��	�~�kr�~�ш������D�6���i�bM%B��@��#E����YW'�����x���]$A���|���Զ[�$4M�̺�j��c%`	��Ӧb&5[q=�܈��!R��!��[����_�,���Y���B���@�QEu]`��l��2��8�m�&�{�US�>�����j�ae��Ff�^�i�_���qL|J�pP�8��i�@�� �œ����R4�~��ŀ_1�"k�f\���E߇A�F!j������|����3�p	GǄ��g4���|�o��������?!j��;c�ފO4�������m6ita���Q��ӕ�<���	`ZE���x-��A��*:y���������_������S\0��K��!��<���Q���c�M��"�'�,�.(�n#d')��T�Y���J����¸�=�����=���s#!w^���D]�,tҌ����܀���n�ri�=�h-�ʨ6��U�z!6�ғ���ٍ�����ȕ�i� ��ʁ���+��=�~��0(�gm��t��AL��ӎ7�7�?m2�e��t�]��q��qE{�	EJl$��Fҁ���uEq�zsM�5̅k�C~���2`^��������i�3m6��w��)�[~d�F;��>��V��Tᶻ��Ac���U��FF֞ڠ��<Q^���k����Y=1c�o�5�+�o���	q:B�˴�gf��d���	�G0q�뵜HT+�t7&c��MIL]����c��M�Hb�H���N��$*��쁻C���G@�V����F&����A��!�F����/\h����I�S:�m���Yg�qj2|�d2�pp�qQb��4����a�I��w����ѥ� �}�W�;�#h���o"u��� �7���f$�$V�U~��C���{-M9�Ƥ4k��� x"�?`P����y�����[��-f�Q]p��n=����Bn� M�0~�W�/��#�qsm�1��'�g.sbK�n�u�jd#Z��
��M�$�b!d��ov��hI�@*�H͡N����v����f���Hh3��YOP-02�jt�M�F�}r�v[��t�35�'��hLS��X���*3<`�����3ҋ��Ireq�ď�2 = �GQpA��ڳ�\����ޯ��z�jP�-N�����_�~���ě�{��t�Ԝ68�Uj����ĭ�|事��K�ep@䘛YO�-J�p������)~�����}���E�����B�����Pc��Ǆ6�BE҅�.�EI�n�������9 oU��l��#g�|�$I/Zh7Vo���J�C�i���<�ú^���Wu��ﴵQA��@�[m�i4��Z8|݂��@!_�˾[�Ryk/���$�b ��#�0��sf�㕻oI�|�=�C2 _n>/�8���t�CCX����uK��"��n'`��j�\��8]��p�<
-���n�7u���xt���^&��{���Jt��m�S/�V���He?i"ޓC��� �zi�9�	�F� ����U7�WW�9)�u�.v:�b$oͯ��6�����}�o��
�iw���z]�y�~?��f��q���
�9���P�
ٸ�"����ō�����@��j�y��w������z�}�D�$���J�q�n1�R�6��V?o�iBU��|�|�z�l�\���>����B{�\����w�%_�E�*f��B�9�n?�F��U�*3#�Z�.���9`_a�u�2%F�}�-�r<k��.e𤪚Lo�|�.�:%v~�)ӝ����}���x�c�k�/����`	�ZG�7N��{�p�����M���k�҂Z#9�$� 8�=���n�ي�J��`]66�	N����/�	�Uyk�7Mi��=R�R��Xc�ݿ��
�v��#e���
}7�5�	�|��b:�nd��-=�^��JU�V �S�ovw%����٘@��A����P����2�(�}N�����7���z�;	���^���s�%g�	���N���Ҙ3��7��ņV�+4,$1�1<D�%a�z٦`Ÿ���[똵��DoX�?r���.���\�%6����m*���K@��E����rfYm�0��C�dhnt�o�DM<���NŘ�	&%��Nu�O_�$�41�'�jμ7m����#1�"%���
& �!�N@��q(S��<R=�ᮙ&[Ep��
�E����,�1F�2J��
�Ǚ#Sy��dٰ�7�PBs�1#�g=
��l���5�>�o.Y7�&s�Gn�<'d,�����e1����NoT����#���#�J�U������i��r���a^�Y4��=�A����%RW��� ,s��0�yB� ���s<S��:�$4~�5��_4�Z�)�Xh���+�Yĵ�,�j��	r�̮�o�`:\yd��Y�]gk����Α$�ݺ��d��"�C��g
���G�R����8^T)%���Y�n�{�$�1����BuA�֗&w="f�|xv+�K�2�\�]�;(gK@�>;�7eIӪG�����3g�L�e�Q0kl�׹����*~����٘����*��I81�N��*+|�}�5 �غMam4�e�d!D�FW;/L��u�)E�^,�%�I���=f#��آ_g=E��mfj��TC5
.����	�<H��e=h�G4��}�|(�����4g-C|)Y���\So}%M#�:6��[�"�9Ls��a�3R@�
�k]��Iϧ���
2Dڡ"1���C�w$˯6`��k뻉�͌Ey	��C����]�<� 2<�s�f��Ş,P8J�S�Z��^
\ˉ��aS!��V�Ҳ��%�-!��$�`����zm߻���/�&<�#���r]yC ~�o���h�����^z[5B������?��h$�)/n��GA����ީ�C�(@�ϐ���|��LJ��?�ʯ&�w�ͺ�������w7���������P����37P�h]��
��>,�)�D
x�|���+�F�F|5z��k��:�x��F�J�`����"��`F8ִ�����οލ���.�wr���Ȟd��g��]�Њޕ�>�L��Ŕ�b�pPԜv�Zy���E����{�"R{GJ�=&[� �90�#?�ܐ�<Ｐ�,�&򊂵(�/�039a���w%��� B���J�m�!Jg��z6��/��)��5I�(y\�)����ƌ��GZC���N����N{%@m�9��B̊�fIT:��c�/��)T�+�Xo��\o����x��ͿA�2%O�D๎
�Ԁ�+�Z�I����s��Q$�+�'31�8���i0��#S�k-_� 6N-(��e�pA=�͹Ћ�n`��\�+����=����DL{n�2�oc�:,�a�WĮ�=�[��69����C�.�5G���~�����u}��ð��_�.�߽�ݲ��t�q�#*����}E{ݣߗ	D�M���.%���H�[�U������WT�V>���0�F���H��
��{p�2�R�o�T���)�GN�Zut]�`�^ifLB֠���~N��,i�d�>&�E�чƕ(|�af��μ�Q0d�aXR,LI8\�KP'����;(�w����E�ϓMX��2N�d:hye�׉��'�w�/��GI.����n{��m;&D1�^�i�ϰ��C��p����(�B��o�N�5T�K�)n��
Wc+��8ש9'kʱ����D�v�_�\�YH��Yd��hOB;|@�K}-�ǝ3(��		�J�4� ٔ�~�E�u����7N0��l��Po7c�����S�����D���h�]�A�[b��H,o��FĴb�%�}T+���F���V|�Vd��X�̸i�2u9��5v���/����>.��偙��&�́tTŉ?��A�np�����d4��-�-F��)k� ��5���2�㱪�wVܜ3(�*�:�O����&nD7Q)͙�X���[Մ�;.�5�D:K���%,<�(d�"�������$��,(��|~��W_��]Aq݈��nI+��eS-7�vdX)��ݑ�1�m���FG��a�����o�a�n(Ov/��6�7.$��k:묑�qT��7�^p>r���'���!�<�P
K�x��e�ke��[4�����@��FL��?bW-$��J�`Qp����e��1�'d%�"J���KA�ɟ����$vC�-v��MK�M�R­d���栺��1���q)vf�/7�[��VW��.�Ȋ��vq9���To�E�6�.[#��̫?ݧ@y4�_��ΕY'�0���&ɻPOx���k�X�36>���9���"�?i������Bx��<��)a�N�}b=����
y|�$nDAk;`@�W@
�Ȟ'. $H�C�N���1�����G�{8a����b6<���so����A��J����$��VWn4�L��B���#Ozƚ��a���a8ե�!N|����q�1ߧ^~� �eސ�iؽQ��5�FW-��M"S�k�H�a_b��=�`��r�<�=:%�^�e����շU��V����.mRL+g�cʝ�C�ge@�p�@���:NʺGF��j����,�S%��2�\�ѫ$��$�E:;;����\px�]�J�%C������FrL�����!Z�V��%�FHHkL�_M��E���'Es
Z;[|�� �$%L�6�Uz�������2�	�.um��n ��X5�&F�ޮ��P����8;}R#��D+_BZv�)�]���pA��Q?B_(����{p-z;��D���Fy�f'�4�}��@�m�Γ������Q�h��-�k��;#�]&'d�g��l��U�5 �V	I퀾��H5���$���ݜ>xg���<��!��/JnJt�V�Yj�C�m
��m套#��Q�t�ʤ4�P��Mj+���BJu������qɰ�ۍ0�C�v�{����W�������Y�G%�e?�_s�Q��I�̂R3`���̂)b$f�v��	e��f+�&?�L����{�l @>`,�P��;�(�*ƾ	}�9A�WgK�H&TX� (d��|��G����`Keɫ��_|�4L{�%�������K$lr�y����{g��^��>Oa%&�R|6GՄ�y;��vj5�L)Gj;/4+��e����{��y����ʛ��y����Cu��K�I[��t��R]'��m�������Ͼ5S��v�W��w:߬�����-�L�5]�	�&L�u"���"�	9V��(����`���Ч�C��O^`�.�2���(J}Ap�U�B߅`w㡻��dA�=/�c�i�V+�ֈMDa?=`�d`�`MR�N���.>O��\)�PΧO�S�y��/u(�!DS�Q�o}�較��F6ɲ��H8u�}�ѝL
/���k�n|�M�����~��
p;Q��U��>��@,ɫ�t�4y��dk���[.
��$�w�e����Wfg�KUײ�+[88jX���T�	�U6��3����g!��s��7�vq���q����m�;Ͱ�	���c��gL	r�As ���L���,��!����)И�༳r�B��4�:�,'��K�x��oZ�d��@'@�$fX2/��y�:��ڷ�-��6xw#�v<��$/��&X�sP�e!�S��eю8K�
��x��ē�<�P�Mu�*����y��?�tv���kGB>��Oس����p`������^=�����ZYZ����T��%t��[��T<?w��jat�r2 ��~|��xY,V"��3�}���¼}�Q��C�{��W�c��Z�<+qDVRX��Wox�5,��D�s���(��s�U��ǽ�q���uY.g\�I�gp*;b�W�U�(X����ʼ��_>>���G��5e>i���_O�!f��xKl���.mp	o|Ѯ�P�Ka�׉�h@#�����'�� ���3ac�k{�yv���k�*K�b����/ ��
£�@�$���8�uA��]h4tP�O��e