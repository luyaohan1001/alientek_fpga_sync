��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���
�yv�X�C��Wg@�	��"�:����"��)L�)�ڄ�5%I���[Bl��?e$skq�͂�Jt��W��״���6�}�p��"[�M����!n,�0�'ɓ����+��ƍ�:�b����)Lw��>��$�#	�xT��O�.���'-vށ��^g�CAپa5O��LO��~$`���g4��<�Z�>$uc�,:w�.?*=.�.c���,9�Ysh_	\��Q��/��8O�j�i�g�Mi�ZVu�������[��@#�!�W�A8h��ك�V2�z��W��lژt�����D�ً����C���:�i�������� 4z��.W��L�),�N䀸�N�e�$���fm�k.��q���a�q����d�뒬�:�	��`;T@���Ʊ@�=��-�XUK,OOM��(���#���ٳ#l?�khg�/iB	\k�M��۾����WF��M�
CH'F������T��O������a"p�I=�)����V���R���N!	�R�1
(���uQ�7�iFS�v�/����?���Ŷ��Gn�J7z%`���s��V����J&��2i8�%1��f{�.C�+H~7����ɱL�5�Ec𨉵�m7yXPܙ�)HZ�N��`�Z}B��L��M�h6@������|u7��^��`��m��F��Fc���Ρ��h�Ѷ���w6+�a{��]�m��ōS��픋���Y��5�\����vRcK��4����B18H���vTg�:5��G6���H�"o�$-��8���0:�6����)=j(}���C:���q3�2)�;��ح���Rx\ ������e��4��9ɔC��oe@I��Ւ?����v�݀�ەYaSt|8JzuV$��qfޜ�3�8����L����b�/�P�Q�.;��W��p��R����Z�/�%艆��Vl��'`����pG�F:f��h�`�dl����	P��A��'�ÃM߈&ɍM���U<��ql� 6<���"~���r��%��K��w�N�.W��y����7���s���3eF�X�H���e��O2|���4��+��Cޔ�������*����F��-�~:jù��x�v���S�<ҤvY�-�[`A�k���
�4�1����\���D3�Q[�vʦ�zܼ���a���`^��� Z?��uG�5'}z�n�@�� #�Y�F�?�U=��%���PM�!'#�����@�)��c�;��<���e\[��T���Y�㌚haB�xdPq5����?XN!�,����i����m��Rw���wceڶ5�����_��,1{	��ٝ��,����}��.�:�\ӑ�D�����a�%F4q��U�K�X�O�Ψ��8Hx/��盩���_8��UѣB|�^3q��P_���ws�a³�����(�R>0�r�xb�yP#ěV�5�)Ț�ۚ3@�����y�Wĭw�4��Bƨ��|9��#&��N������ݬh�[Ҙ[��T<�0K�-��U�T-)U��b�1׫G��_��S��2�pX�]͔��F��V���Z2|iL�_�d�ܜ�����f~����.��M�n��\�s�6x/ X����%՞��@N|8����i���*R�TSqC��i���qE��R�D|�����6e �	Zd�m�ki���!��vm����\p�IG�b�W��b�]�Dj�>��l������v���-r87��F��d
���~4ذ�%ó�P�y�nLۖ�*<[n��);�$��H�7����E\����&)��	'��wD��t��o�`PT4(�N\�=�Y���E3|v�3�M�����WM 	�� �ʕ��/*�st�7�V?��M�9E���t��.�n�Wn#�b��A��N|��sT������D ��]/jP&�OS�+E?���~\��,vA�	�)��]�3���2���?�Z�s!ڤ־�
BgP��~]%7�z7jȱ�`v�;�r��U�$ڐ0���.��e"���ݻ`��1v&�� gQ�������-����`�!�'9�v����+��{Pk��c�(�.̫\��%a�k)�x����|�5���t�YO8KoaA�I޿ô��Sv��VF@"P�X~*6���y��<��4��KG�WKs� ;�;�3�\��\zk�[}?|_: 8�� �A1�Q�݈"�shՑ`��B���=�Q����7�0� T����ߕi=4ޏ��[q ��1��x\o��r���O���![���>�h�9���STy)��2��(.���>�EY�R_:3:��"gu6M���|��M)0s�k�����D��߬�r�k&zy{N%��6�7��P�]�=z?nJ�h4v�]k�g)G�K����E�ɶ���h��P��I���c�8�mxƘ���d=,%o��Q�뗫�X|�}�3"rpvh&��^����Cݗ�#J�Q��
�I�]�Ȼ�w%�i�n�?�1� �C��:z����ᅯlz��ɢ�[�a��gMY?�!��2��GQb��M����ԋ�j�Y��@��v*��<�L��]ڵ��ށ��w�#�h��g���F����VC1-��궬H,�SO�À\6��=D��-*�n��3�@���"�Oc=�/���yEf��[KD^|���X��%9�V!�����2p3�كJuU��MSɒepY�{Lø���՝u��_3\� �4^��0��[݈u(��U}��E?��©.�V:f3� ��j�$�����=��/XK8��t�S�VEl)�"�-�Yȩ9�T�D����>C�>rͼxEJ�'�2���s�)�J�->�R���<��$a�$�����f^ y	̴St.����Q �G;�~hn�g��6�x�)��CZ�6��UbeO 
�>X_�SـO[��S'Z��щ��S��cΖ����NX��|�.-Xܐ羙 �&q�>܆�n�[���$!d�*���Ti�n_��ղ��,�#ص���XV���C�
D�ZW���t:z">�ϫҒ�5��5+Ƹ*_�[jol���S��%Klh���9��a7����:_�3)rض���Ş���{R���!1��(�:���,��ՊJ�mI8N��H�v���[�Y���Xj{]�X��+�/���\�
���Xҥ8��W���=����U��\�R��b�ל���q@�ꥨ��4���C�=�jYTX��¿�iI�� ����On�뜭ڙw�ރ Q�y����P����P�����:U��ҫ�/�/;����t�W�=�]A4]��)���(��Ur�2�w|���
$���p�Xp�5��<�\G���f���:��\wV����5�.\S��]!kQ;�ph�������?%Q\m������oQ0xρ�2��H�^D8y�_>�� �����l�<�tY�cX4������9�X�ű���P8�.�J�� �3*�uQ�Vp���c*K�IaA���[�U���Q��W��sV'b��5���R�/��>�f&_D�|8�8�W�N���=m)��v���s-��A��=��zi���� a�C"ZZ1�}U7)�&s
,*�<J�&�]���gz}m��X��ϒ Wѻqy�'�X?5c� F.���(��eN+�ttw�\C1P;M�Yf�rj��F��y���=�ugb����R\��#�0��}閚�)@+�"�c�����N�j�eg�*���dB�'1T�e���pR�EKY��}����qX��I�M*x�[S�̨�[�����T��a� �X��S|�<����G_"��g��-�K�����f�4�r��O����J��^��n���|tz��F��ya�'P7���*`v�Λ\��E��rb"���c�$L�H���7�/u��?�vv�,'��ݣ}��_H5	=;������a5 ��^���i����S)��]��C$�b~���a�A�n?[|̏dg$�%"�A�r����?c�{cyy���=hO�3U,ͺ$!�ht3�@��_k=ń!7μS�_��5�I�j��G��� �e�BU
#|߽<�%����ao�����c�]��g<X�Q[��T��������#1�#�&���Nb�%W�8^#L7�����p�˷���2�.T���{���g�I��5LN�����&]�]N�r��Ԕ�q��"��c.�<��ĒQ�F�N��/���?��0��,��1��=�ו���_���_9s2R|axy0o��ФH�G�5r0��:o =���ޥ��*�u�w�N���#��dG���#������f���vB���7#��b11�	��?m�Q>z�J{hW���ꘑ>��@��U8�Th	7T�,(��Ցș�SG����J��<f����W*��e��&^�q�e�t7�õp-�?������U%U�[��OOo��Ex��V�#�`���	|�l����w�f���bU}�6��0�T�F�7����7&
8{�0�oTY�I���&W��]�&]'�L:�t�,��ܣ�箳���9a����1�R��b	�A��Wm���͞���HJ�ZMu��i�B.�|w_}��������:Ӭ���H4۠�D?��vq<e�d^R�ƶ���Cu�T�v��qȴ����q���,�f�XdT��*��F�A��
$�4��c+B��"�ր���*�k��?Ρ�����+ɛH�(�E�u���T�(ʹe�^����)!Iǯ&K�t����ԗDtut? /���\��?hV�ɷe��&����?��W�a���Ҹ���L��&�_�E:�p�I��w�C&���*�{Ğ��+a��ų�Yٚ{l�W�(�7y�C2��ˣ�a����!V� �.�m|h���� �G&nm�]�8�G���6�,ol�٢�?�T���p�ml{��>�_1��
�㥥�0pe0Oxz�; !j;"K�yn��V^�2�.��O�}G*�S3��P�僊�YJsϗ
���is���[��4�]T/#ZǼ��w6��9_���s�ߙ��g��5�jQ˩V��$t=�gq�iV�b��q�m��V	6�ɯb��=X$��w�ݯrHG����0j�k��ĳ0{>JV�G��@.��2��+��(�LmC�V�67�Mz��6��X�P>�&;.ͯ#i�D�tݯcZ�h�cT��.�h��,��wN�G�����_,٣��}�8�\�uH��Jo��@�����Q�'Y����vR	|�pM�νK"5��s�D�χO�������^��ᯇ��6���%�d�?��[W�p��@ڪ�" ���d�As�U�>���<t�\b0�$H?�Xb����	j�J�����fA���X�r�����y�����,�"u�d\i��A���f9�k�"�bNB�*�1I���b��ɫ�|S"M7UΚ�1z`sR	��Ʃ핢 �����ϣ�e�����WCu�)�4"���[�,�V&X1X	�K�s&��x}$������|����?�p�׌O�|��K�nK��>$*N���m��x���T����/��j�i��15ޫ�?���:�ɴ�R3/���8{i�ձt��L�ki;W������h�N16%�h�/QqР�!�~�r��G�����ƻ1N4�Om�j�د��T��;�ﰛ��$8A�88�����vVK"��^�_�����;a�e!���G�z�z5֕/`���ܚ�;M��w�?��ѿ��)/�D0��	�����2��p���ܫ5]j��a��"� $�\��z��169E��k#�]�ɚ��;yM?QU|�ab�R���_�zn�~_��ZfmK�۰��;� ����_�/٠&�"1�j��H��Y�.�]�)S�t+�exl�xr
���H��oJ\0����3_nM�P�ȭ�[�̾�w_С84l�	���vCϢ'��<�����Y�o�}C˵������#��m�T�!�̦��C��B�`�ِGn�^�+�枫�b�04��0)�g�ҝ��aup��f��H�J���B{pni�=y��\��j���&�,ϖA\d��5L��&��7!))B���X��&��_޼3��IMB:� U�U��@�`��X\� �xҧ*��8 �mW����]���m����d"�"U��b-��7�(ŭs��^y��2�<��AO������)��O���������;9��VZ��Hz�F�8��U;e��8�ڂ�X�F� �Oa��B=�K�ˍt�C���m�t�=��RPw+�x����e��atR��ݠ��B�w�c������S}�?�\�q�y���'�~ �iЫ7/aP�j�6�%���SL����6#�]t�	H*?��r� i;��K�clT��G��i?i�o�3~����a�\`(�!��O�EV�Y��IФ�j�ŀ���˕g׻�J���@l_��Y*��T��'����l��C!֧GV����9Kمt�ټ�:B4*ę�?���E�6߇
�a���~���'�e���~������AG��?�g[�[�^��獽�
ٴ�5b�ߐ%�DȻ}�^��]y��`qhx�(��Ҹ���"�꯸��Ew��id$Ҥ�B��|���ט�v��#,�����V���`=C��r�*�	�^ȱ�S��\+[��p ��9��v�
Z��O�Kr���lb���$俅�sG4;Y��0�z[f��_j~���4^N-��lR�U���KKyZ���ְQߤ�H(?Urt;�(���ޜ�W��YoՒGqř�!L�Ҵ6c9"�����Ꞑ�GttZ��$�YƳ�EJͨ�N�O	�{?�e��^Y;Y��3f
`'<6�:m랓qk���H��Tg����gcm����8�0z����A�J�����,^���m/gύd͹��!�x b�j ��Q��.�߫�7�v[H����F-�����a+�t����ǭ��(A:�%��������͗iwމ��<b,^%����K�6�$� J�z�������)�;��KYq]�u2����孥y�dZMw�Ęr���q*jy8G=���7��'½vK�F� u��I�t�Y^
�œ_�x�-�t&�������z�CO�Y����W6;��"g������y�	ۊ��7@��{@�K$�E�������`T }��:5�F,�/����|�>QE{ էY �;xe�y��.�m\曂�'5�e\����b`�a���9�ʲ�[�jxa#���!T�D>���o���m�V���m���:�� qy�Gi^�C�f�!��7'�m�b��` �3����YX$��|����_�/=�p�r�}̧���sSjM`l7^����Op��{�k�lX~�#�
ܓ`�Yץ���?k".P�� #���Jx�8ʗ���!GQH��d�2���c�����mݙ$*�L���3��:(N�(8@P�l?�i�#&n�M��8�?���v��-������r��znZ�Z���ʱ��rQ��:��p9����j<Ω�&o>HO��R�L�SW���A	&���ob#Q��t��)c��Y�!<��C��(xu�[�q��M$`��H/�2i���DK�L�m��\�y�S��pRdbXR�2�%�����㰢̉S}Aç��9��@9��H2��q_�5鏬?�.�EG� ���	�C�[�Zڽ������OU;P 4n�_}�+;6��{�,rP
�b�(�#}X[���8��,}��*�������E���%zJ�@'��he7/t�2k��8�QY�8�aw��1x:f�JW��mb).�f)>"���3�j$�5K� }��U U�?���u���Խؕ�&k�>�y�b�Ģ�+�C�$:#L���ߺ�w�i�-2ȗ&�e�߰1���o_4��U��%����a�ڊ��tn����'�J�f^L�YT�����{-~k���9����i��(0}rmQ��_�����<�2�P����x gu4�E�~t�n[��h(0m�:��g
��9�St������i�r�t��睞l� 9��RT�X7��шI��g�&1dޚ˟cOA�ӝ�Fm���U�[�$�������ں��y �5w�q��R�?N_�}Q2*9f8���PE��!��[(+	�hϋ���=�$	��������:�s��A���{5�~�$���w�X��2�X� B��s$�LD���Q���'/zm:�z1�Ü~��Μ��q.$٬s���ݏ�5B�Jv��j6@����;��Z��6�ϒr�Ah�g�q���7����f󵭪��#g!r:Wb� "������I`Q}R�W�sD��N�[�1��;�,V-Y�)�~��G�F�J�~'kˇIuh�����js��fE���O�s��>G[�&������'�s?�Qf9�G��C;2=��zrѻ^~�˯�TJW����	0(�
'QR�"�`*k�E��U��V��ฝ����v���]u�yD퓸��T�B1��(��R��N侅|��'��;5]�<L�f����J��������cX�zdȧC����� ��_���;�Z�ej�����@�@��d�g�[�I��0�w����Nr�we�Ǝ��j5`߄Ra��YP�i�Y�t8S8���W�1���S8g���qM�Ð�K�1����,�7�h�@O�Cz��:JMܢԥjl�T�pTo�
y8�z�����K"�DE����YhU��i��#nа9E�6��n$cW�����wO���O�&���k���Ն�(�5f��}���:@��Z�;$���ي�k��j�Z��+3*���<+��c�'QXY�̉�!����>*�쭋�����F�����!�V�?��OX���̗���Gq��=�o�ŃjKb�N�A� :�l���3��B�uਵf�R��͏��;���<1�t���OhX���3Ɨ�U��1����l�������od��� C�k��k��jTf@�KY�B�ـlֵ}$��T���r��2Sz�̲�Ad^�z��;��I鬉7"�6@��W�o��2̱Z�zyuGe@��@3�Ed�[�i��	�Q�n�3 ���|��fED�s��5WR�#WHM��W�J�8$u���� 8������+ZtR��A���1�e�洖&��]��ާ,T�Հ�iLt_:UCs�e8G+Uw�M����1�S��ـb!���)��29� �4��YJ��0%�=N=��7�0������
�.���}�c���a�
�eY�U�M�ڔ�8β*��g�������p7�]���04w���[��2Dnhk�T�����H@	*��,�@�=hQ��,(���)(8��M�V[z1!�y���כ}d��l����ݐ0�k���!52��롥�L���ol-�<�?�+�H��#^(àڔKgթ�D�\t�Û�^;�](��M�����3I/g���I�H�%��F��&�����8��4}�^��+���r���=���g���ڇ��RED��ŧ�{�P�z=��*�Ћ
{q�n�1�:o���Z�M�N�"����d��@�*Cl��݌�<U�;�dz�ݪ:�v,�MϤ�Vt%3��a��Phk6B�����P�;��Yt�9u�4u����b��r�e! ��������a�K�>	��"�&�����3U�ܲ;���z����Oت<0�Hw��@�� ͨb����EAEk�l)����J�^c�b��Q����ͺU"�3��#�Fb��� �)$4���^�~�,�=�
|e��=%�V�@@��)�^�!L!�_����V��AH��0
��1�ہq�c�� -�-��"�ħH�\��J7'�y>`�y=Qb��,��e�]
�2W���L}�7v�aԉ�]���� [y ���6$/D��Tx��@��y4L�X6/��*�����By>��an+��a_�^��y*��c�vD�`�rĚ`�Ss�_�Y:U� �슛R%l���;U�k�Nhh��4������U��ORÈ�[ z���J�B6�ےw<pd=^V[�W^ՊN����9��ce� Dem���1(ۛƺ��>�	x��,��7���*"s��Dӫ�ɋRA`y��8V�<g��+%\-��"�R15��1�r�`i���ЦJ��⤀�����*�hHؿğ$,#�x��i8ŕ\)-{�7F�\dCZn/N,�#��fx�D	9J��ԏ��bƲ��(�|�Cm��TŘ.�t��3����y�@5-.YϢ����A�엊��1D�0��˪P�I0�1��F�*����E������*-D.��ML�^ ۂV�T�Ҟ�V9��"��{�_7�'Q�m��@�@���4��u��vXBiQ'�zi�
rb��j�0;.���]�9 .l �t����8d�I����p�� R���?]݄�/�R�2����|�5��;-_���>��a�^f��3�y�(���j��5_ׯU��v��w�L�9�ܧ�X��"���S�|v�s��ƅW�U�k/�Dk��X�_�?U�Ȗo�⧅]�>\���I_h染�@+4z�ң�ϰCQG�0������h����L�����>�#�'o�y�^��s6��vG�:s�+aǝ�ut�)I= W����f ]��!
��ĊT���m𮂛��|�I�^C�1�"��+Y!qM��ʵ����lzM[�P�0#'�Œ~irٮ�\��3����S<� #;��$xb��0l���^�O	�@䪃C�{�䲲8z_�|�W�^��h�� ac2�ś����X�Ў�N�ő;~ϛ_&������;�+�\l�qἲZ3���o��r��rxe��}z�[���� M���{��F5?�lb�A��"}�3�1l䛽��c������yF�UdZ��<og�x�>J��dX�(6�	%I�\�t���E���Փ�_y�+Rx�<�U%ER��d�ꃐ5FoJ�x�d���13���4}:%gl�c6{��?����H��0���g���u��f���\xȓ��!)���T����Jm�L%T��	?i,H���&pʎ��h0��Ýt\ 8��n��yOS~O���&TC��xg��xI-/(�O�ͣ��s���^&�T�l���2Kv�~Z��y�B��"�z���n�w�N��f�R�W�����+��j�/�)��
7y�G��}��NP�����ϸ�LK��rm&���NU��UY�'ׁ���خ�-��vN���PT��:��Ҭ��O��&U`��ݰF�W_%|�<T?/�kx�>7�c�kճ_�c�ęͪ�	-Ꞷ�3�������hui˒��5ߘb]Y�����2��FfXW��x0��M���	��S� �De�q�u�KA�;�!X�'�p�9{�������u���\��' ��V�2�cM�>w�H�d�Yԃ_~������w�
i���U�����*!�޼?�����C�yj�"Z�{�zz&��%��1R6��.7�У�wͬ�O�([|����|�>L�W)ѳ���(��5S:��Q4#wC��.ˎ�-����Z�D��p��j�4/חV&�L�,��2���^�� {r�z�SLj���i�$�U��j��ǧ'c�$������8?��S�A�����TA�pְ�9˄�%�-Ag��xG 4�d��
�'4
�jy��Em^�
�́Y2�%_rLhJa�[�5A��y�|��d� ������ᤣ�_h�2�)`R-�R[��F��U�뎓�P�Dc-
�OMՖ@KU������ =w��KG3��g������'�@,tC�  4��, r$�#2HՃ�?g�%XX�QH�x�4� 9(�K,���ҭ'�c
�9��C )�|��˱�wp�j�#[�B��N��Z�A�w�Q^��j�t��T�	���"��ICQ���l�Y�qa7CH)we���7 �5A@�U�\TX����+�~i�y~o�jX/�yp��M��A{��5޽������[8�iUљ|K(��kB��/l���"a� �R�������^��8�8L�陴��x3u��T"���Lam!$�̋le���2 ��������Y��6D���ąn%t�P�������֧+����q��?��D����	�
�"R6C�ș@���]L��ֵ�i�nI�䩤��Z�mW|��Z׵
��4(���}�
q1.y�x�� �o��_��+��1-y��C�L�T�T��OA���U���6k�5�q��+о��.�Љ!��R�-����-�;�zY7�����f�ʁY?{E�q�ׇ-���{�½ëT�t;�_���rj������hJ�)��]Ƿ�7�i�����\]�N��e��N�t�E��#h��5�	쳚���q�#�����Z����x�:�)Ȅj�"��s���K�|	�^>k;��f���t/3׼p硋�o	��M|��x=�7��b�=�w\ꮝT���\�w�J�D�>�w�l������q� ���ZØ2:����BW��HHc̣����6p?x#4�'6V�.,A*ab�Ǯ�hp8���_oUV�}�fq��Y�h����$@�^h�& fI��J�6#h[�X���	3Q�sO[���]N� �n]t[�����Y�ٽ?���zFss��  �Y��$7��ɰ'��ԏc�v���:m��ۚbrtx���^�
��[�/ݍ�;�4*�2�ŏ��ֈ��uvZ��)���n-���L9Oh�������u^� ���կ�;M!�x`k�+<A/����1@,�����p��"GL����fླྀd�`m��Q�W��4�@��Ds�]P^��b0�ʮ�.O��ciY!�ൄ��f�#�Yk#�֜���}�u{DUA�:!��� �2T�}D���.�A�\����:��RXS>�'JZo�1q�N�{�����O����x��Q��`M�N��a���oP�Y�~�>��_	�+95�	�hlN�(�]<UJ�k�̫G�'�VfUq+&�z/>�*[l��w]��%��U��/�-.fS��1��R�F_򇼝� �QY��� p�\
_���b�q3����D��<	�����V�Y��R9��w�Uv�^:��5�[��:g��p���n&����@B�W�����r@��;,���%u�=�M�c�ӰN0VJ?l�U��q`��|E�#���OS@~�AE�� k�(����2s���񇑁�3q���>�3^�Љ>��C��s��|_���Ol�J��c�4�ř:���@�bN�X;�a��T7 �h�g'H
W�+��2�YZ�긊_Zv�2�����,ZB���R�������8@�f��o�����n��ݷE��\L;�^�l�j%�"�m@���>̷GD�`:2_6���A���L>ٙ@;3~���#^�;sL��M"�c�P�Â8�Т��I�#q�i�%d����?O8c��D�&d<����W������|oŏ�hZ��>%�`�b�.&Ao��M��کlۃ�1�b�i	��������_#���c(n�޻@��U���WVa�*�l���$H!]�~��f"(���*�-M�d�p���QƋn�Sr�'�Q~�-6�.��t��W�at	CL�/FS0o�n���W�T�5�_�'�ˣ|�BchE|�'�{uY>�a;Wo@�̬����M�%c^����Q~���O��W	L���/�����~��Ofl���I�GJ�+Oy-��>�H?P��hd��Oa�0�c�>3У�VԀ��谙]��	7t�9q<��q%$��R�AV�`���	��hz;ӟ�lX;	���E�>���@Iڞ��
����c��>�	` ��dB�{�1+�ITX��oo.����#Ud y5!��Ȼ�����0��<[	4||��xi�q����$*'k&:F���üB�D�w� 4Q��|i�9�ð���z��;ڌ5K��t9fQ��T�m�*V �߿��7cmv?��\��Ͷ{��R����)�[/�{%��d7����܇�yFP�(I%�޷M�B�%/�F'{.ɣq���_X��$�Y��?`W�co��M�cM�l=2�M��I��A��vm�.�
/�B�|t��l���`uTO�x,j�f�h�م(��Ga`��+�V<l�s8z� ]�� `pI㑨�6�7�C,:��]^*�j\=��Q�@ӴE��ﬧN��¯�MLK�ٻH#gלGܒ�j��܃��u� �4	�0�(TP�Y�Z�P-;��l��h�0ޢK�Ug��f�P6;7�:��8Zv�?��iq�:X>y��s�E)�)����Q�6���sy�:�T�'�6�������GLcD�I�����|uw�׊\ox�D"2 �.3���e^�xNʰp��ޚ�H�割��CҟM�Q�Н~sd��vi"��N�2'l7"��\���A;@�^��=RB��{O����&G�o+�c��M���-�X��ݷQ? ��Q"���ɒ�/.�b��im	��,Wp͗�U܁W�3��X	��#�B���0�����x��B�"J�V�`u��oe�B�<!�#��`�hԤ�V�N6�~QNM�4�%ߎ���>*��đ�߲�'U��X>�Q,�Z*���	�߀��cf+�]���p<�DE�?1s�m�O��01��)��D���"!?�s�����iTCғ*�;:���lD�)3���c�N��'r_�3�S[ͺ�\s�iZ��yi��� ������"{B���>B;�#�5��eڞ���6�-$P�"��eQC�I%������� H�$V�����_"���ꮷ:	�4��>��M[,�:��G4�OC]��6�{h�5���O�ve��M��}$����6�n��6�Y��av`M9t�	ϒ6��Bt��J3�8�c��_#A�M#m�Q���.%��ב���ƿ�H��}_EJ鯒K�2 � �����;�8�"�Q�Yw��ʝ:�V�Ï�ٲW�10��p��9 V�2�<��J��W��&5<�B���re	,��5Oh��W���t�kxto�O���dρy΂�tV&��ķ&�낷����j��2 �Zᒄ�M�,[�g¤�N�w\�x	��
LV߀ك��(����:�ԿHy�ʗJ�X��)p�;O"�ۦ�V	��nI�;���r�w��Y�_ {�{�|-!%��`�����-j0���銇�;©޾o�/Jv��PQ��+3�.G��-��c
w��g@�>;T��3��^�U���������x�:��pKh���% �r
��S�r4M.��8�������D��!�v�ǝd�A���ޯt�ab�<-�d+�@�f��"��c�f�[�w�|�2�������ߑe����{��2�X�<Nml��;X���b����b?3�������T@�ƿہ�W�0��c
N.
�]��n�;x�u�����ь)}3��%`�
:X��3<GFO�3�֏�j��`?F�0jS�U�C��!8i�p�O��(��^n)�1��1�"��[�\!����i��ǿn�̂�U|?��!zY��EU�!���
�*o����H����z�pW��٤�6�J�4gvÛzkx��W�4Õv�}����v�Z<gۍM.,��$j���~t�2�y�1B<$SŌKY�̰���8��0��M_�جTK}�ΌX�O=Z�[��� ��|鉹N°9�j �<�0Cx���9�6�B�3��k�����g��豷��#�&���MϠ26h�C^hƗ!
����7�x-�(P�ouć;(���� ���c9~>�KG7���i��Wv/!i�|)��L�)=� ����KX�9�YW�%���R	��E�3���t�:������n���P��ݗBEBǱ�T��V��HG|�w�W��iY�ұT��.�>� ��j�6K���?�\�N����r�������Xm����?kHC�bl	���2��Ms�M<a "�0eV柠3$ƈC�B��E�e��r�չ�*_B�?�Ż��Ms�2
�c͚t�W�|h5;̈���W�!�;���Y�D�*J���F��DzD�Q�Pa�\39W�ڍ_+YQ*�4���o������I=�}{�V��}�z�1�6�����lk�_������.L�ҿY��U��E����� �����>��T�ZC�B��a��ќ�M=ڪ���|�'B5l��.���W�y�c��������M�7��ͳh��|8!B��Z�
�_�z��7n&첃�
I���Dk����0X��O�C#��C�{cjkI�w���eEJ�B�!�Nq��?  �w���ߑ�6n�������S��HMDp;�\(&N
�iCD�b�:�m��I+���S�S����a��>ٴ�$}�>��慬?U�����7�c�_����fe<���	gd��"�h��-$�����r��p�
�:\�D+���Y��y�j}JoB�n�{�]�O1�i���mW9*�"�[���"��&��@�q4��%�>��v��v�X0�:���^��r�Z|����<Q�a�z{��mܺ��7#Ԏe��
�[�Jn�ܺa*��r�d��R�G��c��z�����+fU�{�tb�c�7Ę׏��~��A鱮�����d�u��`��lD5B�W�M�X����b\��1\�3����ь~��ԭ�r�*���FBQ,
�뽉�P����*��y#���*�}mX����%���A�I���x�f�g�5���Qf��@j��%��0��{�����U�w~��敞 �)�}��?�_�TP(��E��3�=,N���i艛8�����n���/��F0hb�x�WH�~w$ך &���!D�M�"LA��ϸ3�&���p�+�&���{��hP��5~X��R��!D'��Z�QY�#��	�����^�>����=J�哃��bRW��`��&�a�;YY�P�����.���^ʭ�.�_E8����ć����!�K��������4g�mwQ��/�-��ae&�L	����p$�~�p:u�WG	�N	��跿�1"����?�
�u��҉=�l#�g8?�)�3Tљ_H�{�`��.5O�P���S�����f-.��!B>puu=�WuJx�K��O	�/�G٧�i�8}nN�����M
��@�aj��sr�t�\���Ь�F��a�cλV2(Sc-Gm�yb���Ѫ*���(�E��a�+%��tY�Y�v���,�oc��g�9�6M�F�m$1�[��5����\"]��gV;��s|%&O�6��'/m�����̂3�W��+���s�)��p��El춒v/cE=b����3�z%��W*�d`\����I&=�9W׬]d%����������J�fV���k������	^@��rN�u������߶AW��cZ觴�9�MO��۹؆���; ��]c�lH�&����<�_u�
&J��e���z�J*�^�P�6��9J;VG����w >�@݉��s#����x~D2�H��20�ټ�z�f�S�ny�ܺ��`<�n�a��׎�K�oc�{+Cj�Q������R��k+H�w(~}b�M���/��<�g���R��S��O �f6q�(��x>2�[��VT����U�ߔ>�>�\!�2�_��&�@PK�w��x(nl��I5FV��)��������_�0������-cK�����o�A@��w�ˊKL(%��Β[��rN׵^f�}�VA�G�ϝ^�Ղ�M�N�(B���J��$���Uo�ݦX�\�i�z�~��Iq�@l�p�^G�s6B�g�3(�C�`4_�r�����w��	es>��6��7�s&�����QF���b������DW�UIj���� ��ld	8��(,>:&���r(���ADYx? E�~�����?�gQ��a��`� �ܶ�Y
���$�"?���Z1�[eN�׫ٙ�T�y���R��E���������S�}d� ���3'd�+�6�T��$l!��a�������O��پ�޷t���i�kƎ�\0��ZF��T��k	��B��;6�h=�旼�>hE�Xt�UǦY���������?���8^�b��.+�'֏��k�?�JM��r8,*ʩ�:$�o�
���dtc� s�0+������\ ��EA����"=a�$��Jʺ�6� �B����C�h2���t]��&��m��u=�SB��
���&�(�M�p�hq��ȟ��~�L���Ca���}9��t\�M����y)��9��[5��"�\!{vRMh+'v爌��i�v�I��^M<�7�����1�N����P�*jYZ���y�+�l��$!����^����{��D�w#���D��9[��X[�T �����������(�S���oum �6xӑ#F��l	/�tY�^�5�Ү�9��	����N����G���㊎�*��y5|e���G'D+A�慰+�ZSv���P�#Mtm�7�E����˱�W��n�;��	�W9�7����������2t����Z���{�a�0�pG5(���d�r��]^���
VZ
�)�HNy�!��zl��ո�5��I�Z�ؿ��e"�����o�f��Ɓާ�i��f��˝5�R,Yk"a]$U���Į<��q皽�G��fE�$�TsJ�nm�b��{FH�qN���]�0�Hg8M?(E�7fQ�N��n��%?��K���,+�V�p�lZ���FΓ�
{�Ƥ�Bi-�Tl�,�6�#�b���=���%Ta���?�![�uy}wl$��=����C���F�xru��l�/H���lп�L�;���5O@�IϹ��
��Vu�SZ�h� y�r�Z����N=���*r湕�����𖓻��[ݸ�o;>���Y�kN�G;eEڮ{���4M��M�%$�c��x�o,S%4u{��ߪ�5�D����d�dz�$�ØJW�������Fwp�[�X B�8:���c~Ԩw��{Mkz������oZ��� ��u���ÓZ
Fv��8o� �U�a���{�֩at��Qٕ���J�䱸8���4�j�֑-���)����|]s��
X$��`j�Rt��KRlh���H!|�ئM4�H�"k��`�������ϗ�j
!�[w,�>�d!��8X��af���%�jؠ�
x�����19~6��x��#�m��1�n�w��b��5_����C����¿�^���#lm�s�ZS����9����s�A�m�z��,�?Sa<V��q�)@�����u6'��Q#���m^�`&`s�)ws�^!�<J��RT���B(��߻ޯ���s�Ρa��A����(�@Ƭf�g���?�L��Mw�׊��A;L�0�g�؁�3Y	�{�۷��N_�ܞ�
`E~�H��z�ܤ�h�z� d�o;o{k�a1t�i�V(գC�`��Z�O�Abf��y/み��t)�\$�Q�y���cg_`���v'��¯�������o蕋;�:���H���Iց�j����΅��|��@�l��\j�rT��*gc��ɬY�B�����!P6�fp f��$(�+���k�����M3��wp�ӹ�:�α 4]ݧ�
MB��Y�}Ye'ߕ��b��|A%Y_��rg�8z*o-�@�����V��	�t����c����KޘomC�O�<��{��ܳ�F�ӡk��Gp{�<ݒ���r�|g��]@������Qiy
��vԌ]q��8×B�ӊ��q^��+!i˷��?=��{�Ú�о�O���r��͂z�C����|y��	ͩ�� �U�K�k�����\��?��E;�Y"=�)��+��Y�E�o���ڊ������3W��J	�0�={�������>��jrް۰�dʾ�9G@w/��"$7ltyaV'��gy+!��!���Q��`\2�$Y6�U�kUŒV�?�<�K��7����@u�W�V��9�Z��z�W#2��c��ˬ���3��k�����o�fŒs�D��f�^i��㻦ʺ4��'�y]��G��e��v��,Ԉ��>�" ���1ľ$UK�|Ɣ��<�{y�{�b�s�/ n����:��w�+*~�@Ű����p��ؚ�cY�i�0��L�讅ʶ�Ai��q�e}�f���[D�i�WY�0��?����W���g�(��=OQ���b�7�Ls�����@F�@�r�}l�������%p��Н�T��[W��������5oC=�24":���?2�}�v��ƿ�ʝ��I>�a�u�0��ᓸ0�l#\8S+���L�X5F�
䳔d�E��]��Ǿ���a��+Ø��ƻD����|�"]�_�b����`?7�v��Đ����pφ��?4�&��ت�wp��Щ@nD��x��9^�޹@�� ��__UFڥ�E���0Xl������f=�R�A:��<�^��rPD]��	�t���i���@N���fP�� vI{L����KM��Ē��@u}�߉�j.��jugV�y�;�qmK�X�ʓ%�q����G��P��#	��Wo�z9��,s�gt�;'�a6����0���������1B��$iEd��N�Ϯׯ�gi_a$n�(� Q��cAX��e�]��4�CMt��ޭ<<��7�G��9p+�5w�\lv����3�����_����3(�5cS�߇��[\��G�=�/..�N�k�m�!�
'���cy4�����U%�(�E��7�)q_N�Mk&v��}�d�r�5��,oҦFR�ɵ���'�N��D�x�o!I�Ld
��b��h���$w��y�N���_7���iݢ'+̓�-^��)���Q�L3W'-w��.j4���<�X���E��"�5�����]B�j�%9mn�qgf���>�����+�i���݂�Keq��D�~Uw���drk��dJ�+��\�I�gsH��3������0I�4݀AF�W7��]�o?���Y!5�.�<&̕h�5�=(qM���mu�绬@�T�$����'�?���A��|�[�9���@BY�E��Z�ָ��K�<�(y��h��I�6g�3J��uV�z���1���:�����6R��󽰆�W�g[h�]R���>��r���Mp�
-v�&�H�Z1� ��%	4G��h���Xq��T��.����K�b8��r��1�t��٦s��@s�}Xe��'K�z[36��pՖ�c�v"D���&�����٦�sfo�H^gf�R��W���T�?��8Z+��໡oX�q�+ǿd� o0 x�9��e��%^iD_�,-0y>��>���e~x���
˘��1:]-~��	�\2kmp�]7él*s�ڢ=�6�,�#Ś Ȩ��]��h_�Mw�K���c`�� ��2_Ge�y̓���V\��G�B/��$�u�5�X"�P�F8���d7o�nZa�FB�{>%#u�J�?Ḳ�T����f�d���q��|�����+r�u�����a^�h��=�Q+;v�i��;�k�w/�c�������`f��
\�V��N��C��[�����g<���jV���g�%�ZM��|�0_�i��,h�/�B�~w�}}���UV��e�Q������)��̉`��P��֧��W^@T��D-��囍ۢ���+WYÝx��U}�8��eʩ�C:#w�?O��D� �� �cFB\8�l�2 �F�* ��K�g^rB>Z:�e�@��p���[)Ya�����K:�]x-��	N�k@�V/��T��a^!�y���"7
)|f�>�����WDVt�yY�Ǧ�Rѿ�w��.q����tC�l!�b�����=�\�� &N��`C�#7�h.�+>K�;�qt�,���SCo��C�W��3~�d�1>|O�|�oᘀ�\ Gn�*~/�ՙ�{Z>�@�� ��XGMgU9��vgIirC���&��