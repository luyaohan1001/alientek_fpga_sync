��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O����<r��[y�$��l�`���+�=��/9P&�~���ƽ�������3K��=ˀ �I�?}��@�_��-�	Q5v�M�6e>Tţ����S�俈��ևi#��:@���u���1(�����]Cg&��iAW�9-�;	0n|��������ʾ�E����l�*_��M���hm4@��mP�h?ƩRyj��;�ְ��������= /�T�T���7J�c��r�`2���᎜�8m�X]�M��~�%F�h�|�����6�DPy-Ɖ����=ў7r[�	A� Q�N�2o�Yx��g!B�g��N$��#���56amˉj@��QA~([��/��N�]���D,��	��I!���G� =s!���oܪ!Ȑ���y�&��8��
ZH�������.ua4��3-RNN�iHD�F�W�$g%�i�T?͏s<h@�����^?	��%���r@Oikc'����j0Ɯ6k}%z�A9g.�e�N(���KZu*$DY�0W��p�AL��P�^�eDZAe����f }���T�Y�o�ĺ�耖�e;�]�l�;�n���a�L�P�$)���O�����5|{-m��D�(�4��P{��%���Q¬'',P�0�R��q"w�44,��
A�P�'{��J��=��Rg�i%�z��]˼���&X-sP(@!;I+t%�N�
��eG� t� )C�H
�OJT@"SXV[H��Q&��'�KVw�N�w���>�L��:$B����Ǥ\�\�q�\��J�t����\�5��n�5j�iiq��+E��(�sSH\��W4��l�/��D�O߇T��xR�
��=�G�������em��i~�4U:BX]S|��S��!���M�Sr�M_��&�⌑^���p�_�Wm��*�t���S	 S2��bO��n�n8@�����m�1��2���պ4H8�u����XZ�Yt�w��Cuy#����HA�I,RH� ���"�S����	�-
z��T��?qq l��f�"��q*!�6]�s��ɪ�[��<|M6~�n�P��bM`�ibUB0����9�C]�dB`���s�H+6V!�ƍTo8�,Z��>@㾐� uq�2Dh�6#f���H�]j���R[���&�.'�V����\�M&�������Z�Bh�����cJ�z���<�7��	FQr,;��*��,i�8�pt�C�_㶬5��X߉'��8�Tye��Ϫ�W���+f�-1�|tHu���*�K��)��8�E ���x�eEY(�_c����W7�X/�2N� p�[���� ��*��Qxϩ�Ae��L�bg��P#�#�GM�SV_���uK�t���Y	|�W�dc��ɯP�����ihJ)a�FK�DD�h�{���cA�@�<����;1@U�k	���7���\�`��^5��"�b��$q ZՏ_���h,8oF¦޼�dh3��Y�i�.`Z4*���O3��m�㇉�R�	���ٳ8T�x�¨�T��i9,�ʂ�$<�&0�:\
� �p�?�%�T+�$��1A9/�?Bz\��aA��cE4QZ��FF2���s�W�v+�؈�ઓU�Nr��������@t�B3Қ[M[��/@Q���pCoP��4����$�p�T�==�N��z$;��"\�AJW�oR��mbd5��q����I����5�Kh�QLq�� a�o�#u�t)w�C�<���wqk��#���U��x�KDd���Q�� ��k9����^d=��ս9G>x-�7�s�|(��]��5C�(���q:>;�I�\0���YYt�����:2)�d��ɋ��1�kl��j��,�bDv����jH3��/��z `[�ײV>ti�A�u.�5,'�����:ߒ3��q_Y�{~����-M��rvE�n��6	ld�G)0�Li����+3��Hp�]^����Ab�![���y$�#��]4/V���L�G�m�0���ۙ�eD�}6�ݛ-�b���(5!n$Zf��͌�:(2�:�s�i�~3���fx����)_�J����w!�qB��"|H�����q���������p��"��J�}Z��S��V�����l\�8贿I���ۻ�? 0A˥ȁ�8�t��.97�lr~�՞���6�Qgt����A����Ѧ@���`Ax��m���9�	oz`�<�E$��ִ�&j�ð���5��
V�Te�?�g��:��t��g�p2ԻJb�!r�DC�}��V]N�}��ί��d��	ŕHq�z��}@����#�t��l�HK����E��w��� U�!�'W�َ�h!���8a�Om���9���3a�����B`f��h�Ŷؽ^����6��N����U�Sq$l�eI�u�L۬�h�~O���̙�i��)��Kg�?sU�Y�"�-/�4��_m߂j�E�>�d+�x�����((��%M���x\v����f>�^wH�tw�B"�T�0	��v0(����A���ᖆd'e��F���¸~�H��2}ED�~�n�L�3n�>m�l+O�۬O�W�1�j������!O8�!М��t|y�I4P�I��C����p��X�4^�|���0l..xnv@dq���*����6F����{��گk&p�եL�f�P�0��q��!�Nȁ����J��`b��R�4���\�7�S��G�/�,�z.������~"�I��b
��A$�&f��xP%��u�"t�\ENm\[q��J�m�YX�Lw[HSP���|,��y[z��L�D2�?K*�]@\dR
�p�wI[*ؕ;%�������n�L*��(Y�T0[�[�e�opu4�҃�pWɔ���e�F�Ո[D���ݖ��Z9�����p��侣Q�Cj�E�������9��FF��x1c~�C������3J�N��+ ���"�7�V�ѱI4�kQ���ʃ�Q�j�V_�'��T�pʷ�փuI���vw��E�¡�����J���7����������?�XC�����..��L�
�\>�Z#G���a~k{{5닷z�A˯���萹��XBj|�`��
�\�<&
�9;�(�� �˃�8hj��l�'�]�W�,��&kz6�����0���e[��������
ߎ0�Y�s6W�Ğ�^v7�(x�%�P�!��g�z3g�Q��Z|+�D����~y|fV�&��L�q�Ȣ9M?��R([u� ߳V��CɄ�`�¯��uRZ����v�u 8���`�d�t�`ҁUu�\+:�D����|�p�| N�����jpU�;(4�kR�drh��4�8���ܹ�
�[�Ј�t���KD���i�X�wg ײCd��%l�,�1��c��9�,Y��'r�-���u�?,��!�)���H1~��"�-P�&��,��" �#s�����:"c�~Ƭ�k$>}Mڎ}=�,��_kYmE��IyOP<F�mR7�1|IUA����MY�d@�ۋɧ�a���^���]w�����!'X�oɖ��Oi`��=u�۫V2�>)i��<�y���q:�.�jM�ܼ4	c�$E� �˴o"�ǝh�.�Us@EM��.�TM`^W u���'ȴ��]�*��|s�D������s�㟈������Z�Lׇ|�W1�2p�N �?�%;�K�?m�5��T�ZY�j���g\~�l;N��c�f���&nb�Xvīxz^�RZ�p|�9�7��O�@������l>3�OZg����,x�'f�/�qe���` d"N7���B�*y�8���8�O]I_@��j'֔C�w�5~ �{�'U�la�Ր1U,m�g�m�L��	�4�C��R�c�O�X#6�"��K�@:6�ϽO�x�Ē�?]>F9�"3�r�2��λ�м"m;!v�|,(x0�^����f��k��k~�o��b��6&_�N�|u�ڇKOA��7�$��g�?��M.ar�)�w��g��rO�<��_�P�'�ϥ��N��%T�����r�,�ih�U�6a��?w��3ԥa�g̙[Z��O���Л���M@s�K �B�[���9js]oYj|��<	��
M�Β��|"vU^��֏�wp����2_��<���|p�N�����WϞ��ʦ03LmI�2�@H���y��A���@٦��!6N&����E���נa)���7�]�����*>�.5h-{(����T�?pi����қiN�jW�V����A��B��Kа69�1Hg��~��b���˂�#���p�!��*]�Wk�2��c���q�����*�q��R�"����h�e����d��
�.���W����t�` f���ڊB*�� �hy�e���Y�l7L�.qF�o�P�k�Y�se��
s���B0����r]܆�iƁ�]�&!���Jă�nHb�&���0i�̈dh��r�}~�N� �7���-	^t�����p������㨢N��c��Us�L��˷6XH�?�I���tF�}
:oh���+&��z�B�si9z���Df��'O�
8�z3�_*���'�o�2ܹ�2�UI'�o��ԧ"*���� V"�n����H��./U�-m�����@x�-y��s!H���a��(���]���h���Z5���	;n2��K�{^Z�E�$���3qT��x�����Ok:��v��;mwd�FQ4��uk[3|�S-������g�=�NƆ׺E� ��˵��Ͷ��������	q�9��]Vbgx��I�b�: *�6WQ9���D��!���g�^��v�2�I��@�_*	�bX�9H���u;5k�@����n�X������g*�	�-�t4��R�ƪ�A�<��>�2�%4�e=S{�Q J:���D��]���qP,�'�.A���vj���}�WF_�b���ƨE%��Q+�������7�i�7Q��Jj��VZ�����Fy�	o�<��s�͸{�� ��4�3v��ߟ
�D@!<5o񆙾�E�Q�[��O�i��ِ�4PW�*:~��Y����h�y8���'/��q����(��/p,EM%�NB�賑�>6)��1�l��Pb�� |~kvw ���ȿ�]M�ٝ�@(��u�ʳ�l��n.�"�ƃ@g�A>�L�)��N"-��2�\�-P&#�&W�Ua��>D[8�������D�����,���cSŧ)2�=*����2��mAug��rEr�F���C�9C��"��S�dA�^�o��{]C��Z�Q>p� R�h߱f��0��W8��ֿ"���.h+V7��Rh�bx�Ů͔r#=+���.�K~%c9���L��D*�)_�┆���̫|z�������X���qm���Y�͙�W�I'b?"���_4������&�Y��K�氷����D��_��%<���2#��\_UzP������}n=��+�%:3����0�� ���;ຈz�v�ӭ&M���f��B�T���_�X}�V	��[rL�y+��=��r��
{���|�ތ�4� ֥�2�O���7o��`�~�6�{���[�X]΋���_9͂ZU\c�gƚ��q&t2�dX�c�������ǃ���i�2S;�Z�D��=��j�E/�x뼪�x89�B�fE�
�[� ��r��y�s1p���π���Kڟ���1&����GC�EO��ATW��Fr�����N/���J=���u�,MJ���W��X'Z��(�H$5�.�n�"�j�5�xmN?��j�6��O�yZ�����揤�L��1�'Ӿ�u_�p��E�*��/�޹oD��_�5��ӻ���#t�	�)L��)pI�;���ۋ8ѐ��&��['*��E�ܔ�إ�(3��b���������J)�P
�S�T#D -�������˞:���#?R��~�Rj�4��꬜�p�3� _���B�y쥛�|ʭ��=�&B����sT�fBg6i�[�-��)����LL�x���$?�N�	jh����O�	��W��)���(���<ȸS�\~Sᱜ�`�:���e�hk��3��Dh����y��R���v"w� ����E*����œ:+�{�U�-����L�>��������&J�2G��ju�MP��*pY��z���v��2�{*5p9�������[�¥�-pmn�'�����ڡ�}��BGRdt�o��<�Al�;���M߅�hʲA=�Ta�PñyM��m4[z�K�0\�TC�x��{�������h����������S-��}��1����WO�O3��W/hI�����.�
�
9�
�xo�z�"��D�*��.�4��?{:6�Pg�K�iZ�� � :�_�}���D�yzhq ��%�47�`L�Mc�@�g���z��S�>7#�ɓOa�����09��D��m���|]�{��R����}䔕p��/��L���n��y�#��_���QD�� 1Бt�P���TS�l��퐒d&nc����2�lO���t�h���p2r?�U�0�g��~r5O��.�TDhS��	��$�;è�%8��ݝ������F�d�,��G�6��>AM+jG�q���:as(eW-O����hfUJ#���8ԗ��Hn�U�g����G̼�͕!-��l;�Ƿo=���|��N�Nf�U1S�W�'�C��H��J�/�<����heKn�vu�R���� ��;��>Bi�|��"be�����6��:�g�Z04s��/�a�;۬���d|�k^8!�aO[��"cnz\?��W
Y��� ��ky��2y5̥��o���l�` �"N�rq��f�(�� �_W�Q_��"���v����x]�y`&zkL�A�@3F��M�t� ���T�cҽ?7�d��$�V��רGp�E����m�2����7�<��G���/�x{�L��͌<�E)����"'Q�	�S�H^_К��w�e;�`3�]�<C�I`Ʌ�rU]�ݸ,V�cw�L�i~�U[��g�}a��}����^Q�n�ݥ�����O������!Nwa�oa�`0�0�I���$�mJ�C1���O�4����m[[c�I�WCa�&X)g������"��J��I�Tc)���U�����4P� �u��f�%;��8!�+��mG�P��YU�A��cU����ګ�#��p�f,�^v`�=����)�wc�|��L�DY\i;�#n�B�Xz�:[�3�37z��g.���[�\��t���G����{�;�����C���c@H��c^X�J�	:�2�ʣ��ӵ��&�����*�
Gd�%��ݍ�}����ҟU�Su��D�A�$��|?o(�F��|���.�j����f�������$gˏ���T�͋�7�A��&%o�~��fU���X��M/��4�Dt9aA�i���=( |�UT��
��pB��e��I��;,R�����I~%���8@�U?���_�9.�zQ�*;v4 ��5-�����r�>(�o�Q%UMk�6�#�<��S���W<�3�
P� �(k;:�X��	Fw�H$Ǥ�8U�,Y�Y\;�ҭNqbl簉`L�[/��L���K÷�&��xO��j��R�;���Ⱥ�E�xf���f[K�)���Ŕn���})�D[0?���`�$���i%�pb��
z���7�bj+f���FyAEr�d�c0vYa�@�4����m>�O
a�/z;��r�OX
���w�iv��4H��+�^jɜ2>�o���v,�R��%��������T�:�tx���Q�2_���]7^����ɚ�e�~V�F𯨭i?���}kY� _��A�+02dr�H�@�N��y���_S$�A.�Fg�83���l��v�	�l��ٴk����������{9������
Bۤ�$�$>3�;w '����3Y?�ᛋ�Jg$��!F5s@��^U]�P.�Q���p�2*R�cD���*e�F��6��[a�0�qd����꽗��vrO���N���xS��_�7{��/9D�%ur��u��n�a�7�Yů���-�Mc,�D熒}�*^�R����[� 6�iv$���	�O3\Q�_1Pw�(�����&�'����	I�= ��H�'?�z��p��099�HM��;�;��CB.+o���LpL%;��WB��R ��o�������Q=K�ƹ!�%[����ze­R6qJ�s�ܷ�PEtǹ�K9?�'M3��e��=�����+��l��D��7V�B��ݠ��S'0���\�a��6�Q*bA��iB�S����#|,dm������4�Q���6D~Va��-���9x�9���D��ӹ�`G��V���r����ؙ��fХM�Dr�T%���X�Nˡ^H��q� @Vf����Ȍs��(�>�rW����곬?��L�J�p:]G\\�?׋J������莅^��w�x����1�p8�A��
�����p`���zn�b��E�����vui��غ�;���f�D�+�O@@�P���Lf�8Zö����
��3bx�	=��aH��e��T'K�&�����pH͙��|ީ}[]ם���I&�[�l�ȶU����@ƻK^e
Ǫ�n"��>蘀�[E�.oH��jl��֧�,��1�$��@m�~a�=�gP����iy�>�N�+��rT���Ca|G�\7�UY`ح�*ԕ8�Jj�;ˠe[�nH��0yy�]-
<�g��Pb�ec���cү	�a�i��Qe9FR&��rq��ߞ���4��8�v��Ţ�m�vP��
M�M�V���	ͬ��x�������;B�Nq3V&%���d}tKs4�<X_%L����AK8M?i[H���9"^Z� ��x�MV�%)h�>�D�5�Rb߂0�MD�]�l��x�v�|���"�~!�bn��f6������Rsņ5.$�Q]5UsO��6�Y�֞"�A*�6̮y)3���3�"��y�Ƶ���Y��Q쿢%�f9�s�O�3��~-YUэ�֏���.((�G��E�2P����i�oʫ�Ѡ�X��oՆ�/̰�s�4��s��ujh	K���u|Cڰ`�]T���^�<N`ӣ�*ۥ�(8j���=�8z�~Z��/Ҕ.�h�e��g�m_�Y���=�Z0����H,Wa�IiG�m��RN�m��S]���ҳ���>z�ǻ�~����rE.��|��r�{�3�g�S�e2��`B�ʭkS�#b'z����Z'�u�)f�բ7�TM���R�е�k'�#�=�}	8�hHa��]���>�n�����zb��MT��f`M��TY�~0L\e�4d���<��G�PQ�
��-�n��T�lg�hF[!-�����z�T�D�-p��}R	�����S�wϮ�� �z���V��N�fj.��{nZ��G�^7��	��m�P6cמ
�q��4n�f7���MT������"�0����	����7���>H�RX��bT%��I]o��!������c��|��2_�K��b K>���-��=s+ҫ��Lz�.����=�y4EO[�m�NR����C�	��U������I��}*��&�9@q�	5,\/����"샊��вԵ�
�B�3���q�T��g��⬴�[N(ZZe�����qgף���l�?�q+>���B5��^FF��ٕ����kHW���	A�r�ȁl�^��r-n�i�N��'��q\�bS lَ���i�auV`�wdBR��"$�����L'9��OU��Ɉe�R��ӹF�=4E,�	���	�;d�!>�z�����>B�0���lW�ܽ�d�گ٧4��cm����+ݐ�a��R���V�>��7�o.�?ˍ�tk�<G8-��q������;��8���@��$��UH��Шl�s҄W|,�T ~p3���S�A�L���;����ADSRxF���5��4�9=w��/�;�#����͌0�� /�
<�i)Id��f��v��N��q�A"�C��>^��ThI���d�ej��U�ff�c�/F���s-ه0��$��#�_���[�ވ��<�D�F>"/�A�BE��YX�v��Lf��*P��Qo�*�e���y��xc����s��,xE�	������(��X004N�Bݙ絞��Ln-�1�X�+���F�­�A�I��f��,�Pi��W�@-����!��)�.�Ѧ��lL=����C�(`�}X���H�c��r�Y�'_��� �垈U�{׸3.e�l����"�B�r'�d����v��aa�)�M/��1���E2OI������볲�F��#i�e9���'Z��C�u/n,HpW+���I_voXa��$��i���_ধ����Q����Y�qd�m��������Ɨ!3����˶��+P(Ŗ�Q7�,����8��A5[�%V�����ZZ�Gz��(R����
�X�����;�:W\�qѥď�yfa�(]��b�ȼ�Jڝ:Y���`���3�c����g�ZI��UO��FH=ߍ����}��� X��o�r>�E,��{����B�-����^��>�v��d��(,�=����w���H�~t��z�*ĭdj���vԐ��V���V��\��-��b.�潍� �0\ߦ��P�Z�^�^b��Q��5��R��C	�h�x�?�t�����B���/̆�]Ů2ւ{ь2&a�S"���0p;�h�'l���B�U�y�@HZ4ja)1�Bܮj�2�5��0K�o���E�ƞ��i�iC�MF��� �:���)'�"G^�z	t-%~��#B�zV7]����̄H:���<L���U訮3��<]�绾KD�J��5�����(������2��3id���L�<��
;H|w��f�8�[�/~�w:��?]ĉU�>���Ed�̈́�0�0ܐ��J��#���u q�1�q�ߓ��AQ�ɏM������ؔ_'�W��݇A��z�tq�,N���R�a~C��m�(U�_\�|��M��N!��"J�	�{�f�:P�k�[ӱ|;�.��$ī��Pv��I��z{�`E@���;{����k>#��)|!.��e[�	�W���<8l��O��M�d,��6K�^�jM^���9j�MNQ��Z�������:�w�8��SY����>!�p�3V,��!pOBT��(�s��V���3�6φm�p�aI^
d>��r����pfs���dϊ���d��H��R�
%okL|�Rz�/����e�r6�@��}<H�Y��
Y���c��+U&��T�yS�!��	N��w�Q��Ws��
3K�4�UD����k5���6���cf��y��2���Z�1���yIT�!�r��RܸՔ��hʰ��昜�2F�u��7��]g�J�����E_W������o5C�~��ڤ��Y�$��aď<{i�IK�����N'�B�P��n~ys�CMD��bY�5A���=�$��'���׷ٿ^�?�7��*c�|yIĴ��|nD�A�ψ}%Ļxì�q��R�r
���0?T\���OA���4����p7N*���Oͯ�9pݽ�4�E����J\���s���#�#�ʈj�01}ҥ��b���<�7��zE�.�+W��
�M����"����,)�j��=��� �h�㽑pEE��������n'��(�az �۽�c�h�E*}Ep)����ST@ЁMc�������⠝��#�9�'wio.�)�@��w�-�lU־*���d��y�[��?�>�6��q�Tg 8���N|���N>���������m2T�b�c�k�A0�.e���i�g;{�_�߉K놞wm��He������*�߸D�����"�P�G��_\*\�KUp�#��H�n<l	@cQ�B@��R���N���޿�O�n,���:��C��)� (���ª���@:�ld����u�n'�X��Ǔ�1�A��N����M�i����r�0�v�۱�m�Ku�i�`/)���U0m�`3~wG<`���,��'�:��|��\
q*~�֑z����8�_�G6��.`)�tP���r�G��檅��E�Q,j��;D�����k$�С�Ƨ��T��?��
������J5�~�#��s���ϑ��x1��<e�Ʒؤ�跾�K���`es��4>��!9�
�o���G�-�4֚�lP����◥�ȋ�'?Ϙ��#�sª��fu v��0�WI�b�7�tӂ�u�4��^����R(��nc��:�
��z�ƯUS;�( ����F�6z�V#@�M՛��r��IsX�<gS�����jZ_��&���/Ϲ]/��(H8Y�}��w�v�K?�xY�`�������F�7A�h�+�a��}c�X]-��0���f&��ZΉ�"3ģ!(���S��"UiM$\�c�&�=R����*���QQ����5�(�QA̔�Z%C�S��Hh��G�#�ʲ9r_��i��?}�s]>5c���kc�6�zI���lW���S�~Y�~)�
�t,�����9^�������\�t��w�wb�u�7*�3�t��s�Ңj˓c8[G�(O�qv̵5���s:������+��NfC��L� !�hw�=�[�z�}�o�tΰ�|�dP�J0EJ�l�| ���Q����0���d8���E�@�4d#��.��R���k ��'��L�<kd�����%|
}�SŰB/F�i���B�瞧��!�z\׎�V�s���
�*�XH��3�2`k�Y�e��/�
IwLNʶ����-e.�5��MmF��jȱ$��!հ����X�;	;?zG榀y�B^6\�A7��*k�w�35�́�,V�)~����e���0�ƴ��V����eM��z ��{����
�l��;�J�'\a��'F�`}Ba��ݖ��5�����{l��h��H�m��Qh���;�@6k�Ϣ�bKO �8�:Z��^�V��S�n� ]#��.{�`�&�E�2�||�J� Zx��%A�t_�ȫ37"$hXJ���z%6���K�ԩyzF��-o��S{��L�\�\�	�H��BR�L;����Ii~,7uy�o�_{q��\��M�Lv*Qq��жJzhBK015��,Ͻ����������rc?�.��W%f�O!��Ź��Lܣ�E�*�,g?�1/��̘�i,u9���l� ����;���9d3-�����9��6��qO(5���+����yd���^75�ګ{��R��틖e	�s������BO�Xّ-~x��J���uq}�鎺����z66��;W
7�o9ǥ�b��ܿ���c:\�+魲�	�p	ķ�0-=�����<	�KQZC�J����nL���-��2K�}c�����%�s�޸�0�-.T_E��UV��?)w.����&�\�`e�ݑI�����1��@|�`��ox�'�9X���|rQ���f�VW���>k��wm�h��;�*���g�JФԖP�L.ݤ��a�N�m�8����������Fs�� �݋idf�+�8�!�;�T�O�Ý��4��]�=��hZ��׎:�-w/Į֍mm�A��Em����(qH|��'\����c����ߊ�B�nn��Z��=��|�B����u�T�<�H�A�8�X
I{I�i����*G�y��2��k�LKUl!�ͫ����4u*ƭ��qZԼ�����Jb���pq�����R3*�̪3 m��fLr֦0qK$�"!Cg�Ԁm١@��'�IcȻ1��q}Z��߅�|���gc�i���\�lJH@���f��=����������_4j���f�o>��9/��IR,Q�Z�C<Y[�������m��v@#�u,g!���nW�;4*�ܤ��x�/X��d��6�0�!�d-ҥ�g�'f<��:j4�8@�YE8�y�L���;5�Fo�{��I	� �O���?F)i���wo��/�S�I)͵H��\��f#�HFɎ�j���z$�V�fv��XrcW�� *��'��ae�B��cG5` GV����t"�R��aկ������HuH���I$=����ߪ��������Ɲި�w��XFѩ�=:�uv���Ls���[Yf�!����X�zco�i��Ym�U�VG���I��"5�{n���
�,P%�/1"�հ��w c��xSx�w�R�r��3�v�&D"OIII�-cP�+k�o2�~����\j�Y�� ?�dd�W��!�]��ӗ��}λ��_&�A�&x��|-�Z���-g�ɢڪ�
��t�����Fa��}�f}6ѱdFȯ\V�>�!���-�ѯ�B�;�D"g/u�4?#a�/B(�t��,���Z�
1�e�������;��1�W��Z���;�)W�.͹I������z���/	B�PK�� ��'�&qc�-�x���1�mI$�ci%"�;y+;"K�CG���H�f���x����c�d6�
h��C3ae�� ����1�#�su�5$��V��;��RY�ϭ)@����\�~ޭ���W�:�Ϳ����`,���ysX�·���Üv�غ���7�Ji�E�*c)>q�x��/;��mN^�=_�ܑ~kh۳�ßY_Ț�hx_����8����� E�;:���>��Y<"�'_��J�adt}��D�B�h�C���l��(${\��4��m���'iI��d��V���Nċ��򋪠E!����2���+�&f~+�Ը��ߴ��*��xS���*F�3tHM5o~|���
��Y%�V����ٯ
��;�]��c�����1���߇�M�!&�{xn�NN(W��,�����.�Ҧٮԓ��6�ulK���BJ���%�b�L�P�7
.E	E�,Ԏ�˅��;rR6��S4�����jD������anH�;4���z����.��2���.Bb�#� S5s�c1��
������p�$J_�p�{q(*��:�/�RϢҠ2���@o7Y�I�@�rl�"�
��S����������LD�>l���jDk&9�@���3cu��<'�wo��qp��d����4\�
04�n�����u!uؘ�a'�9�D&��t�)����P���]>a$f�>�36�A�v2�%�*N�7��/,n��Z�cM^�nS?c�M�n��X�hD�h8.��|���>u��o����de^Co?�_Kn*�܊Oޅ�O�����X��[�x�Saբ��������0�SA��h�$��\%1o9��/�he^�(+��f3/�9 }^�[�hi�̾9����5���йχ���Ir ��f��C�^�������|�	(���7PŬ_�ݸ��m�[��Vc���[�-:#X횙���<<��X>�:������`��Jb�O���7��B�ʯ�^N�� ���c3�F��*M˃{蒼4sQQר�"j�����A
�t�,A2��Ⱡ�V�EU����|��՗�ja���'Ց@����=4j�)�M:1�J�ǜ�&ߎ㸡֝uC[F��kh��uF�H�i�˒E5�4!?B��9×B���S�ɋ'�"�^U�@\�Z*1�䌵��{���*U�~�>�̢m�'��v@:�%�ʇ����f�~����j��i�^���+�Խ�'O������Ҕڌ	�^
�γIU��Puc�-��9��I�-ɸ������{��a���֭���f�c�ɡ䔖}8�ᦿ,X/Q' x����}4CԖ�q4��<�ۋ���=O��i�EG�I��T��U����qh`��ԍs2(�o��hP�K������*��S��������81��a�D}���h��P��~>_�������_�/�]�k�!a�D9$OI����Z|+Н��>M>�e����m
�FC�@u=\�Nm7�(����Z@i�7���1��=}��d8�Y�\mە������<ʲ�����,1�D��B�.f���S�ƸH���pa���޼�r�~މ����~:h�Z'����j�j�0�Ņ�L	5��dBp�`��]��D>g��?��\���e�^Ӹ��#'�����*5�L�y�	�b�����C^����
n
 �b�H#��@��9�uW�����j�o�I�9"|�׭�P�]�v�,Q5T+ٵE\��bIDn�M�+��1��=D1\��4�5�Q��8��j�cH&o�a�dI����!AY�+�����7�R�C@���)��4s��-���I�=,c��e��w�p{΅45�nJ��� �VQ���:K��@� ���R� ߓ*@q��ּ����f�����<y��xS����g�O��׏~}#�qs˝���8UN�\���wQ���_��Y�p�f���z�>]C�ˆ=�}�ȏ}�-� �f��DG�I��(��+��r!uOd/���ǪqYq��j8_�Ӊ�� ~�<��l�W̤^ޏ�^����m�%3�b#:�X܆&�+5=d�9|R:7N�iT�Y�L.�+1]�K��0��T,z�3=�dp�b!jKj�wk:���9ų�%ROǉ�Пr��}�j�>��,��ޡE���{�r�������-�W�Y�E�����a�Ep��<1۳y��$��
r�/Ɖ�m=�68�Yi�ߙ��>�c)�T_���"��W�	�z6\�;��W���J�ld1������.��^Jgr�\�A��{�x���	º���=ί�E��Ům�k�b�6l�0�������L"������X�ٹ�v<�Ls=,���}LgZ�����J�
*1N�M��Ձٌ�y7��y@>-M�⤨��}�GW'0��6�_��{%[[���#:�6l
���o�S� h���vF�p(ܥ���P��ni����u�k�]|��٥_T���/j-iMM�g���s�Nx-B�i���T��p&�0�alt��^<�_����>l�C����f�G}�<��^1���[�&�уg~���~��� P0c��;�C��Y[���C�V�Ƒ���k��������s�,��K,���m��g�l� �Q���;��c~���T��e�E�0�z�`��_�i�я!���>�"���v� l`7�[�W�M�Us��1=��+� �4�&���������vdv��ݺ. 8��N���9vӂh7nW�
���y?�2�����V�$����}�s����Vh�~�]���%�@�*G����[.d7��|���R��3�W=��cv� ��:H�<q4u��C����8sdZ��2hD?�J8��Mz(2��i����H hu�hʕ�x��*
���a�95?%�M�.JT��Q�BFP0�>,3[�j�����P�$S\Q�r�r�QV�v8ɺ�Bi� �&�$����q5ˈ�x1AC���������
hȬ�9I5#>��q�C#px3�g�<�-覸����uH�����K�g��P��c0bN�����cl�Ѫ�j�b��qA���8/҆��)�uo�]Z�Q#/BY\�uGˑ��/ˈC�u�x�Uxn��8-e�Ü���~dC�ґ��/E���e��y�w&2�'j��N;�n
�/�H#P!���lZ����=B�{d�@��	�=hg�K"�c�#�~�w=�Ќoz��J���#����R�o���%�*,_� L��WC�,���ɟ��bɤ~��<��x �ƲV��ؖ[�A����'��{��E���(�8������w#Z�R�Ş�<#G�x�j�>iF���L���
��R��0��R�Rv��C��X���8�k)���6&!&}xdx�����4?�Q�5	jU&$�l
v���g���앁����YJ��Iz��\�D�Smm�%�fJ�-���_��B�ȣ�СE۝��ħ��=ɩ1塲�G��gÄ��&2��n�Its���ԪFF*\	lX�r��5G4&������}pe0/�=s�����6Û_�H��,�B�	�F~n%�B?���8㝆�>ޢ���&����Y�V;8�4�W0x	���~����-�7�l�Lo6�F5�#�@�L5b@[�v4��u��;��x��(>����p���2ٲ�^�|�BD���8-ՙsX��7l�BFz��cXY�tIJ}�wI�lu�����pk؂t�7:f/c����u�T��������NEH�=k�l)a&�Mz+#uL���O���$�9�	g��Hae��)�05�jؘu��Cߓ>�7SdEݥ��H��G�y"��|�=�o�!�����Q���qK���9)>\ݍ���P�	��o8��m0���c���A�� 
Xs�YZ��[��^��.�Jo�켍��_:�\���,푟F�ڂqJjR̵-��%hG���g�":>�����L�u�(�� ��v#�0���D�9e}A�Yq1�ڙ��e��"/B���:��m��A����դ�:����'�ǒ�����,?���X����wҐ{4��K�^����u6��(��ln��.F��1��4�aJ� ���>.���=f0�Z�DZ��|M:�4�+�0Bg3�'���sJ��U��7P9K�R�|/��Y^�v"hc��ɱ�BP�G�1�&"��vP*��9�S��pp濼�b�^;��QAͼ�c�_V\���h����U�j�[�����й^���i%LLH����3�J��-=���N�o�%�.�S���ob� 2ʉ���0�z�v�	�e-(�u6�\L1[���%em��?$a�P|cc�'޼��	�$� &`�}9����Z˘��E�1�+���mt��yIM�����_Ԙ���+��P���9�WK��X��x�d�bq���ʤ��}���r�(�r�4�!u�)t�B���k.A+�Zݕ�t�|�$�^/w�誉H�K�1Ӷ�T��?�4*�QS�#:TM�r�����ᵃPE��VZ���-RCލ�,�.�d�����?|轛挹퐘}����;_Jǳ$�##���N0��]�_F��<�X3Pi�������$��p�E �P���$ڻU��	ƪ�
:�H�by�t�3E��VοAH�dY���<"�7��g
B�cP��p&�����3#/�J��Ka�!���pV��7"x��`,�uH�s�Vt��.�[��&g��څ���]"6P��h����n��!�(�&���^B����շlE yC��s��(�#�, �>>���؜��i
�xǱ+3���D��'�\�W�����'|c?d2���#R�e#u��	��7�E�h���75j��Wx�,������H秲Q6-=Ɖ���Qn_7����`˃b}Jԙ�Ӽ���GB�9����OXXDy�,�sɥ̌ļ���:���v��K��'�~��^]�:{�����z����{(�����ѵ�x,��'��b�vC�7!5�Ai+b��ȡ
G���M�}��1C��k�� eQ�t���Z��R��0Xɰ�V�H0��L�.{�����M��� �J����}z �2�{ï�JN����=���.;�p��J��청���#8�76t���Έ�և�%k�T	a�#��1�ө=ͱ_=6�M����э��c�pE)7���D��\1+d�.B�� �6��һ�^Z!��*/��	!�;���c>r��Y;��'<R�[�Xk(ǯ]���_<E�@N�C�wL�Cz�%M�}F=�+�k��P�k�Ij�������?�S��[1�k�8wb�ۍ����V�ҲZ�)��G�y�5�`�8��c��Ͷ��Ð\$ޔNcc�x:~Q�qz%1;´˕�Xs���z��~���񍶁��̷~I�b��o'/�O��k��<#�R��?F��f����O%��KM���N����ػ*�0��`W�V+W6��b�e���L:`�#���Y�MC! sy`�lo~��3Z�� ���n�����z��i(��U�?�?a��Cb�����ߐ4�0��	XC+u��];��fS{(��r$�7������FC\�>M�_As�OklUY�[��y&`�S�����.6��"�߇��J�B",d�@s���y��3pw
��I���GR<��<Ⰰ���b62��_Q4�}d<���n�*����W�I/�q8��ZGb��,�]&�U(%^�9�L_�۠|Vf����	�cҢsùOP(��
��j�hfui>����MS�u��G@�S�������ݏb�nFv;��1�� =W�⽶e��}N��w:�=v5�pN�t��%*8��ɍ��W�<���O}�JS��3�MnP��3P;gDn ��}yz�}G���og㴄 �j����\�;�JJW����G��OEp��ʪ��ئ�M� �o��$��x���\_+��Td/W�A�����d���2��a��GfvJ���>���J,Y����(�=���w,�.5ښ��:���҉�:,"n��z�][�$�m�p1U������2��IX(s��ȡ�?��W�����2g5 �j��V���Lu䭲xi�1��1o*���O���k����P���}[���x���J��P��]D����L�L�V�B�������Q�42�N��d�CI|�����gäiV�Gf-G� �a��7���0�5޽����KB��O��Jo�)/1�oy�����h�8���*�%���ҵ02,�,�V�N�k�*	��P����A�=���}s8���ƭ����6�v�O������b�������&�n�hZ6��P��L��r��:0�~_��-d+�6��˞���w��h�{-rEP���v�8��q�Q�5O�;���{���b���4�������-\����2�!8�w�v�lb�h�y�2i��uō��Ts��a�����H����i�\��
n�:����Ko,���C�-Ub�5e��+��e[HNK�5KQv��y���4��ps�>i9��W�R��u!;����8Ն��[C��d����7��''��-�5Zw�{/��E�j�͋�K�6�HpG��d�<�:�7��6M���!�靦�������G�U2�v�����uc�%�J)�=��p�L�L��&��tapIS��6�>,��]ʺ5�C�v���/G?ES
�Evf��I���8?�ȇA�b	wXNt�t�g����C��>�D��v���u��5��M����6��Cu��&iVPU�r|��ة�9��Nu���	�;�&!Ei�)Ti�(:��,F�qzd�F8��e��6d?�Kl[�,��;J��a\�^����_�IbYTԛ'k��W,6z�����IY!�I��4�;tA\/q�TO�����8�y�x&�����un�;܏^A?�4IQ�%��g�����9�&���(�(��5���QvY-e��Q9�Yp�p��p��xL��� P-`�uS.K�Ee��k1�8�^"V����~�"�Wk���xÝ�����aT@�]��L%�%i4�w�D�F���)��_Uog��v�q*,��/˩	�1YH�IP1T�̆z�O�˺R'�äͽF���C��0��}�4�O�<͍��θb���.y=�'�O�Fwm�=T[as�F�y˟��?I�J6�NkBx��V)�6�����@Rz���:H��?҃b	G�'�ӽ"��Z	/��${w*�~o��>t"�lr��#;h�^���j�N7��LA�	{�g�C�sl��I��z*{/��������d����EB�{l�}M l����\�1��;q5l3��5{sj O���m��"����q�}���*�>u*��gR��5{��{[u-��*9.�N�~F`�ꦿ�/�D����ך��k�D��]��"�:����Ѭ<"�<Rd3w�6�ۡv���D[���$_�:A"�H�j#m�����P��#Z��o� nQ�*֩Xζ�N�gLV�O�b�O6�d�D���̣�o̝�|mRR*АL\�%"`������o�9* ��V��R��6�g��@bg�C1���w{<�9�;+;[��hn�
�+~�
�+�B���������>^
`;0�E.���(��o�^��-�k�~[XA4rE�v�zqH�_����ڠ�m��d�i*U�
u��2������0��D�>ڷ:�D�2����L<�k��`P��^�n=��E���D���kM��ᬵ���vBV�R$�Lz��n��N֟a'��g�K�%iLJ@��e�s������ծ�C�ZVE5�CIkb�oL�t�D��&})d��u��E�+����`�]��:��?c��3����p��e���%
V���fy���Hs���7��v��9J���9b��f`���� ���C}��:��Z*�zf�:���<��?�1� ��{�U7K\��u[��(�z�6ɅJg��1��� �����F�D��k�l5�M?LyʺC\r�d�8o��f�k�}��N�_B�-�OL�^��x����=���U�n�1���䮨����ЙΥ��1i�Ԗ�93���E��,pՏ����O�)��vr��V�y, �f������6���EQ�v��G�<` �3rL��<Ϩ���M�p��A6�Y�D���Z��1Ǆ��F	Z���֬�w�B������ ���ƽ�*{m�t�u
b�d�����:h�ga�/<�������	�����䅺(��X�������J�t�1Y���ۮ��W�gg��+��m�z�
��/!��"�Q	�F"��U�-G꼼^F��/�������Z��8r�_D��S�46L��ݸ�D�^܋nw"1׾)"k\��/�� �`�@��5��ڸP=a�%�N�z-��K8�li��j��|�^9�9�u6;����|.�;ڊb�?-���CXm���B\$U�L�gŶ](�{
l�^�r�Gq��$e1�XQ-��gL�W=;%+"(��q��&vtɽ������ǁb|��nN���=2:�o��15�x��������ztl�a�*F��J� R|��=rڽ;�(4c�\����n xNO�o`�����7$q ��q�!O�7��ӳ��S�?�.��)��$�pqOuO�%�K،z��\&��̓�%�<M@����Z2�1���R�����7�D��73H���/�B�FѪ������M�cC7�X{GJ������g��PDF ���	(0�}:t�*`�e����f���H�ڣ����Rw"�����I~��P�}f\�G�3H#	J۷�{��>��6�
X�����}N�\��P������{���q~��3o�.,.�kk��q��~�v^�����[-a�>�of�����[��mRD���i��{�4*��9M�ۡR�� f�?BIԭ���YB	��$������ʔ�'	��b5fN��W�S�d��Bk�hjE������/D�U:��<����R�������IK~�v��k���o��q\$���M��ރi�h]��f;g�^���M�`E�1�Y��<$Kf�� �Z`:�Is���\d��A�WM��3�o�@P�k#D*��#c�w�f��������Q�4ʗ��SQF&.�z��h���o	8���l�.7[�Ao�㛃"���&�T�&���%�y��cm�g�'���(i�%]�z���y;W<W;���g$�v?�����[�/8�m����K{�̸��&�M��:�g׎	4�҄T��fEfgj
��o8tm���5�9��K�
6�+�4;O̖l���}�W�WȺ|^�`A�W��Ȧ��Z)߇����S���E��,�&�
���+L�	�_�L��ɰ��*��~�:,[��ؠ��1��\��������#=Z����R5�� �F�&�khg?6��Đ���M��-�����;�pv����U 8����?�VgO�̓e������m�O�Ra��x=K�m|�����ڟ�y�X��S�M���N�l��{.�,�p�'�WҺq{h��0�s��~�|a z���N���84ӒX���J޴�[��ZS /�I��7R�����\[��5 ���9}򁾖=k��m�I�k[cm�%�r�Wq3��P��t�*�Y�!`mX=9����N)K�]�!K���-y�}�Y$x�&sw�j
��wH{c�U���>'86t<��0w�a���pH���E�%v�%��SO�0�X�C�cv�_��X��qN�7�\�@�v��f)�[���Ҷ��9�'Nن[P�A��=1��P���[�;�F(g�x���ź���"+��s�2��Rt"74�� ��؆d��'I�>�/��^�������k-��zZ�?�dU��v�^6��Xi���bz\5��=�=ة�0��+��{���ә��NI60֤g3-��s\�E;�e.��sD��B��(��~%�_�Ib3���r�~8F2��c��#+�>O�[�c�2z���P�{/���Ր^Ùa�o^��Cg�dOq������qF}������\Zȣ[�E����@�O��4�]v��D�)U6����Ve�$~�c_���	����^K�y�aLֈ��e\�$��h���ۼ/'`\��V�Ѳ��ȒM{���
���㗣{��aDy�o$H&�u�?Hhj��x��jَ\�u�������TX��7�]�t�]��Qj�{Q�ꥉ�	nfw�'�?�����.�(x�\��M>��fl(&	��D��F��gT7^t��;E��P���}PW��<�������.;7ҍ����S	hr��ף2[5a?����uU�������+�N�w���[���i~?Н����y��g��`��KuJH$��v����\'Z�PhZ,��&�y�K���@a����~"E�=�o�&��A��ӏA4YGи�h�E��G�T�������H��5v�1D��&b�������V���Xe�*p����T�X�V���Iډ��%�V�ղ����������P�v��0�O��K'�֤n)���F4�o�!p��R�$�vv�W�T!��
��v8������j.1��o9	�I���̇����ZCmvP�P�4�J�GW�<�!} Y�\V�>y���#�/�6F~���hD;A�U �+��1М��+s_�X:{�c����ظ�Y��C~��� �"��ud��q�7�ʤ9u���T�չ8!�}�5w�52
���<�>��:���a���f�[ow�}�g���:�n�S��R��mE=�)�D��]���<�	B�M�Z�F;5��Wn��Y��ZTG�?B�P\P��fqV�J;�aQ�"hڳ��G'XQPƮxlV�Mq���]�s=6I��h�a;��"� Ef�Q�)�����Q��Z�0_0�,�Dy�Uv��e�a^�1�W�iN���l�$d��g���U�[���wM����J�`���G/yfg+�/�֦�E��U�ڂ[5���qu���u^-��q׭�	��U�_�k�ٷUlEe���s����v�$ ��-�i��k�Ÿ�?&��<5���Y����=|�1��.L;�
<}�������N��pyd���T�=~��Td�T
��h��i�!1��s�>����z[�ߏ䱉�Qb@�bU���PJ���,۲1��{܍��d5ZW��KG[lQ�IK "�y�9t��0>�ll��Lt���y������9���Γi�G�z=�j}�+hkAK�kv���>���E�IK�6#7�p
ݽ�h�!g�
��y\t�ɌŦo���g5:�g����Q����D}mhM0��yZ�cKSi�ސK�jy�a��'F�d���~;BO��h!Nw�̃��@<���L��l"��<L��=�+�Vd��g��}����|��*1�m�V+��L/�y#��_�fD��*Kp�9s0�^�{o��	�3:y������"���'����,j6�}N��O���ᛣ��D{A���?�B��J�=籧E�`>{�����ԫ� W�D��G0�.o�=R\X-vD
�������:Wi`K��ܽ���|�"�A �]-di}/���v邸���I+���Hx�i�B)Ӳ5<�SH���s�NN��'���U�l���CeoL�IA��6b�30�¸p}��(H�B�D:�с�&��ң��ɭ6��!=�	���� l�'���AD��n%+�S=����<� r���)��홲v��㠄&~���4T���z��)[jM�I�]���j�S�K�v�*`
�d�N��x��Hf�	��O�T�5�A�/�$JX��cۿ%�!���cZBcK0��j9��R��˜G��DVJl�J����h�aU\��ϖZ}���KT�wD�8\:���0::���$��Mu�fc�L����F�bh���7��wB��tz`J��-֥��L`�Q��ʦ�p��s=_�{L��:V=:��?�WcX����Nk�Eα�e9hlމ�����b�^C()q�i�H�0����eDVF�7nsn�j����4g)�X �V�LtG8<�I�IT�Z���z[`n��ҹ���;k�]�.�
�M{���-V�2��H&�ǁ�۹rR[���'�H�]?S:�$��r�*�}�����w�s�ȵ����~�� ��P��!<^��_r�qcw�a�v?� bt��@;���H @�F&##��z �4���������W�wC�&�6�~�ݫ�����+�_�RʲқW�-M$ȩ���Hۥdx`�E�]��#>-z�� lL�/⎥԰�]Ռe�N#��K��"VJ�8�����C��1�-b���o*`�&���3"?�z�
N�E-#�38��
�)��)�w�XP���t�[��y�1MH�5֊��6�r�X�"TY�2}7�C�ɍ,[�-l�j*�m�����p�<�e@&}�d!�2K���=�E���"�q.��Eܚ��'B� ��x���R�Q��9�d��E�1�=Q3v`���o���y�o����D��3Iu�`�Ԡ~�pB�ݑ�LC���-�0ʎK^�ԟ{���>�Lp�,�r�H�Z+��`�pc���b�ߌ��;�Hj�m�v��T#�����@@��(����E��������t�X�2�q��<�L��!u~�>)抂�qR�A��<ca�)���a��H�/sW�M����|-�1oh���*��"-}a3PhH�.�oL���]ߩޠ򳁿BM���@���/���;k�������3���ج�Uķ#E�ahHüz���j�p8�*dw��G<�!Ca�5WA�U�x$*�ص-ʆ�*�B1�'A����-�������@�C��B�o9����Q�n]jPw�Ђ���n��~�aj@�P�}f�����xd}q��C��e�o��x+�6!M3���=�������q��\.�J��	(�aHgJ?^�ܷ��$�fjh��Lu�N���2�� ں�+$��_ˈ#��:���3�Qε�|��|��;D'�M�/B�K#/U���'{rSt��O�{q~���-��Dun����e���IeDI��{��ڌ��vd��S^�����;$U��>�1�r�W�	L�6�8et���a�4H%���DB^��*�zlJ��~�� ��;ͽ����ޔ����w�D��e5__v
*y0���=�brt�E�����L%\u�d�Q�2�o���-��}/��W`WY�.W��m=�/�p��ڔ��i�Ga���[��m�Bh5���,G���h������W�CfxDσ�&�A&��v,�)��:�IDe�8�.Ԛ����1/�ay/�=]�w�#jĠ?�D�|#뺙	��HH)Ù1_��n΢H��$�k��wW��l�Ϛ��N}IC�V(~A�[�)Ӂ0�:�@��oa�U�aNݕ|!^JӘ���B�� ��cӂkEbF�@d�t��BY5k���䕅�ul��ވjjbw���d�nB�8��WC:(��I�K�����RH���p��,�.YN�s�z�a&�~��	���7Y��_l Z%b����MaV�#G��:��J�����BV���-�kA���l���Q�m8�`�.GcKeb6��_fb4��Fo�)�A+�1s1!�Ǯb�
����?'Rj���s6Y�W�_�P���1/�����N���yI��M�6M|��x�S�2q��������"�	8+p@����5B^>�dL-m)��!kG���W3��}��N
�s��CzǊw��������ɴ�Jy��C$��|�5a��F����Τ���!�cD�OKB�bR��JUsˋV�:�������r�Ӄ[xԅ3n4��h=_�9�'fd��[CU/��,��Ce��M��.�8t���d�M}�w��]}TO�����T<b�v�q���3wp�]�A^ Y��Mԅ`���6eC&;E�n�~�nt`�r]�]�����p{�/��k
��Z�����09�����_�q}E�cw�'�+�U�{8d�]x����ty����q���]}���Ag�3γ�`y2����?�����
��]08����8�<C���'�5@zm��&ɭ�c^�c��9!E$�N���t����Q)�����)�����$HW�Ӑ��8��Iv�Cp��Q�x�⣊F4�o?C����B�Oe��)P���E�9)�S�R�׆�-H�O�k>|�ޤ�jiM�M�xV�^:�K�(�Qn�L�h���=�r�H��<F`l�U���j,��	�L�o][F2ϭ�=,�����v��2շ1ŭڌe�L�U߮���A�Ui��������0�ϳ^�4��;���!^�6��R90��:������/�9jH���iC��H�=����Ν��O�%���$}3N{�S����/5�n���0X� :(r8_GNNԂjJ��h���N�}u��ș\���͵����@?۵�
�/L#(���&�Lu;��pn#'jUlfho�Ʊ��8��>�O�	vi�܀4��=��qf)5f;��˦�U���+���;�a1X+E�f���6Bغ�#9j><���Ҷ�0-�+�?e�-5�ct�ՖB�ƸE�}���y�x�G��$F:Hے�Z�+��2�Hi%*�ٖP�SyE:6�߻��㒧w�J��`��c�"'���|���S� ��s�Un���$O ޘf3�x֏�PPeD+��[k-i��ZL+��*g(|Z�n������"Roe�o��{��8��w|��Ԧڌ9�"�P�hKmU�-*
�-K�1�������� <_?�F���q���ŵ������T�L��h���L<tV����ʑ�U§���k(�`�8K�*m�ǿ����)@N2�VW|v����;GC�e�����v�j�DF÷��=��s�1U���P�loO�I#�bWO�3�j�� ��W��%Z��E�j+=*& ÚF�����#��N_a�?\�Ŵ� ����`. *%�!`�9-�'���̒Re�֏8�����V�����|��K_(�?�����G����[���{^%�������V��+����M�9�n�j�!��J��lu�<5���ߪ�i�(y����E�֩�	����g�z���Үrx��n%8�
 �;�boN��y���pI��&����v0��:Ż�3�%��Y����~�`��Z����*�q�i�� u��Ҽ8�XPiG`�$�AN�Y	�Y��eP\��Po([���Z$9�S�Ŕ���u��R��Z���z�4��}rsr���ݜ7���p�a����;�6�
.H�t�e�*&�i��7Zk�̽9{�0�{׊�Zַ��N#pg9S]w�%�g=�5�����C�*�\�#s{M��&l��+�Ծ�l��*�#6߳G�"�J�h^{&
mO�K$P4�M�逾�D�h$\]��j�$:�}rW��nTտ �7��"G<�mB�����ý\|��k�-瘔[W7�91*	0�v���m�N��sC4��2>BЎ��8��)q $�+����/�&V�/~����+�*y�A@|�~�k�&�O�1jo�CH�|����w�j&��0:�.?*B��N �mL�ط�D]�2ь��o���Q�$�D��@R'k�m�-r�%��3�<۱���R�]52`�ߕj��'P1߫LG8A,�A�J;�:�R7Ͷ6f/(��'=8D���)����B�.��e��3���<���,�"�9ѵ3�A����v`�g�̥�[�q��Vp��౛5@���S�g�Ed�J�ge 2���@ځ��-7/��*���"�=r�Kd&Q �՚�f��UH�B	�uR��rY�ڶ��U�~ N&m�y�km/l��\���q����a��fq*'0�,
�SȢG�y�+B�2��,[��Б����w�7��/��gA�����:�!M�g��%��gZ���Y��s���p���--��ۆ^Κ$9񧷿�^g�[*1�'���_������:'b�~����G��M�P�@�R���-=Wh�u>}��;��t�ַ��cf�������߸��}���He�S�i���.}�6�C�Č�w*Q>(�7�ƏT������8Y��ʳ�рPt���Y\31��L4�������-|�l;�Z��V���|m�<�C�9t�L|3�7U�ϕ���$*G��%��N3�Z1�B@�pC�f�{4��!h;}�~�m�}ѹ��钔x"��}�/ �À���k�����&�&�/�8�^3U*!��Ǹ��3���V��m�q�So��dl�p�����Ĭ�U͗��$����N����#�[������P���F�f��x�I��ӷSQ@6ܔ�A�,6t,wG����6���ȿGT{Օi�����N �&@��qrx2cr���_e��J���eC�H޺~-�T4����;Nlθ��!b\>#<#a�P�I���H�Az*֞�5XI��8�$k������U�=J8U�=CDB���w�������{Oa\C�G�:}�!�F޸Z#`O��M��K�L%�"��W��.F�I���P>��g��YI�J%0:�:̴r�wـ |(�Xp���Yro��r}S�P��BE�	v�-8��x .Ls�6g�9#��	���Qh��up��e�%���O:@��P�n! ��g��>6�ϟ:?}D�S�Q&.(�����C�A�˚��F&�J�CM�]��c�~ ����W�ZU9�3��m�X+p���`�]ֽ���ʔQ_Z�-@qVCն�	��d2���<q�9J�P�F--ā�k)�̻\�F� �e��t@�ө%���3���r
�u9*l�<��؊u�JWMٟD��p���n��Z
w���~=9���,�mn�"K�@+ץ�KM�D������	-;.mT��U�(6�I�V������L�\�m-�.���h~��(]ŋ[ਖom5�hs,��+f�@�ݭmN
K@;U��g ~U��ģ�A]m�T��>ƌ�x�|M�T��D;�hk1dw�R�&�b���	�4�zԥ���|�ns �G��#�W�Rm�I�E��a�=�ؙ���r�����B�G��x�$��3𕦯�s��_)V��s^ϫ/����m.�J�0�4���{r���M��kحa/�hT�F�e�Ά��ݝt�p/����O�$�IS��,�/p1���`��D������O"��6�:H<���0'�Z]��驊"wS�j�rq���\r� Q��{C%�%#�"�������Y.4�1�іQ�l��^�ʰY(�t���Ӓ���<�a�b!J�����}��o�>���1p��	��T�E���:�@�$)=ڤ��x&hH �%�!��|Č�v�HZ��f̹�6�=��h��,>��Rg,�������<Ln���|Q�+��s���%$U������\�?�����$���������-:�F_��KLT�2���>yk�o̩����Kl��ht0��?�
��t\k�Y��^�金(�u7�Q��g��x�����O���wa��cז(m\�/~����ک�>wcE~J��#BJ��Ѫ�x�7.9�x/v��d]A<����t��|L]DX�xW�#�<zV�]KC7�AO�q���M�f��w����<�u��34&�Xǰ]J.1�qVLn��
��nteۤ�ed�y�6�F�G��M�D�"��R�6��I�d���6��m%���虖Ż$��Ԝ>�e1����z�W��M�������-Ң��3'ܡ�/7E��WR�~��J�p�ۺl�?�
�W�/��w�@M��t�7?�_w��[2<��,Z�I��e�'�,�Ӂ��Rg�Kp%w�����G���'1��EK���	������ ɛdE=�!	��?�Y*���P��h�N~ۀ�Fi�#�X"�h֯�D3����ƠW.��������r���d;(����ٳnc;��>�'26�˨��)�m�����S!,ߩR�r�N����!�CƈlQ1q��jZ&�?�8"�d-�
�O;Sk��+��EX;��sjR���m��Qpz�t��9O �0�VQ)�Z��$��4��=o}�&M�ʓ��ٿz&�h'��o�jV��=�ՓϺ`���1�YH5��}à�5��w�ʛ��&=h��u��V�h]�����ZΔ�/�H�qn jA��i[��T7���(����c�^���[�a��nD�t��� �̀����_�N���]Pu�8����Q,@ie�>F��w�K��LzҨ����5�%L�Ӂ/�������i_���m�+)΋��J�5�/��	������������kJ�������נ��]�7��Rp��oʩ����+|�Ȍp�
,<�Vn�ȹ;-(]-迱,��+Xxʆ����� Ыna� �p-�ӽ�{���$D��nqlW+���������璢^[DB�g�$@���T5q�����\�#~K_�O����Eߖ�ۍ0HEl&�o�����qG8l�F>�P?a1.��Q��<��("�؂�xӌ�5�B���tr|�bZ�����p��[����b��E��W:���`r~Z���)���Ǣ,��)%�,�������8b�đ\���b�&jl۩�>S�!,����o6��>��l��x�|�Z,�r�;{��c��H��Rv�[J�U��GG.��feˣ���8k;�aX{Yx>��c�lI��(c��r���T�A�]!���yK`4�$���%*�!O���x�;��̣��3��e+�fmV&F̯X~���r'χou�E�+3���Ty��2�qR{v� [x�8s��^Pu�>�95��Q��'��U>X���x�QM�v�������U��|�üIU���o�	�q|��%DR	����ᵓz�8�����iՉ��1'H�&���|ࡿD��6���`�G%&��K$�l�sJ�m�I�^^�3AkFj���K����@5X�Q�K�x��X�v:(�vܹ�R�Q��оQ�2kj;ZrC��Μ@�λ�ҵ�����9�B�$ ��.^Q]V/�9�h������E��ٝ�s�'�Y�&���094�&ϳBI�*Ԗ� -7l\��oš���۔���"����hyj̐;�~鄞���Z�wf��Y�s���]??�m,��	���@�L"��,�����i����:U�3�9���C��u{+d�P������&�"Uz �-NPV:֐�)1�0z����]��SV�����[��|ʋ�h�jx>ǥ����=�m'k�N(Ps��K��� 29'�6���fm�S�Qo��Z�8V'؈�}Y�i:��E�1r��7�3r��yt���0`]:�'�5��yiQݞ�J�n�Ou�t��:����#s�mEJrn�޲�L�ͭ��^��SW�3gk�
hw�?�0�reH���O����c<����<��6L[�_G/[�J�`���n�$R�N��6��v�G��gdZ���q�F�����gXn����0���j!�A��C�{U`�2�iJ����H�8�9�<qbi}|�Gu4�Ұ2/�%~hz'Ԁ��6)Mb���b
��ة �y�1~���>�� ����.R_M��6$��'��vVz���L��tUx�qq�#�sUԿ���Gk�2$6E��4+Rʥ<�����Jc,�N��7Lj��\g	-.{F�%>��V��2��5�8���E#9>�����G�Z߅pn���̌\(��vA^,MO�o��
~��~U�^-0�wm��K65��?\C���(0���5�4Dd63��ګ�l?n,=ΐ��&ӨJ��1X�Es��,���mS2�
=;ϯ���i��q+ޏ�Q=g���Y�\�Y�λ,��B+`�$�����¥���;�wE]���@w,fޢ⠤.�?����{�M� w����W��Ez*� q^�`z�_��G��:�u_�-p:
	��Ù�V�rY��!A��'H��m��U����T�8�w�%���cK]�5r�b�ݚ�����e���� �z���]��'��c	s',Q�E�(�i�d��Z�Bɽ��.܎�E6�T��G���? y�l�ʪ���0B��C�1���E��<���KO�G�N�'�c��c����0�e5:Tm���l8B<F�	p��T����XE��aØ��*Y�?_���0d1����X,Xă�O�P9�/ÂI2^�*�p8J5+��\3��F�T�˚����b�(�6\@Eo"�[�����}�=�3X������ʺ	��ͬ�И6�S�"�:;y'�mQ��9o�H���^��x�dtB�s�Qt���]t�*0���ڥ�=F|mS�Ӣ��
o��o5�r���C�@��cP� *C���p�)W
�PmK�Rpl-(�Z�7 �Z~4�Z���K�x#z�s�d�b������B+�R�:œi[o�P���/y^��b��{6u;|�����"l���F�R�P�0XK�_��mհQ8��`}$���eeD��Z5�Nz��i�����)1)�1���*�#��Z����F�R�^.yJظz�>�"� �{�N�k��y�mn(�|lY`r/t��D�3�A�{B��=>M�{*����N��� ]�P������kx��20j�����4�n���>"H�ޙGUh����jW:o�?5����h�_��d�< D~�Gk�����C��g�8�(�����H�[h�r3�a>�,�\_w� ���ד��썌r?�R7t�n�i#�~�U-鵙���T�s��p��9��E 7�x�u�pҋ,U��T�R����l�G+��c?�\7�����~7R�T�1�WL��D��/͈�@�2P6�6o%���f[H9.��=��O*\��>L6��0ҩ$ga�{�}�?���\�� �o��a	�	a|_Fʀ��}��Zr�̅-��ذ{l',��'��`��N�9|JK���l[�A�kJ���������: ��<��B���f��}TZm+�=kQ��ӢS6:��mS,u��,CT�^ݯ����m�O�7}�eb�(����!I�L��ЇS%Y�J�$�
�X"Wv�j�_B�5|\�
5�ٜK�A;A���H��%�wOa��<�CF�1#����?o٬�?����V��$�_IE��;0 �Ъ�a|�-�WL��TUu� N�ot�$ywo��Gѩf��~m5@�Ǩ����iw��?�K]����a�x�?
��Z����?��n%�Z���:��'�xB���ƭ��G�G:M��Zc����I(����6c)6ˌ������/�g�F+8x�������|Yjm���ˢ� �PBe�x/,OLjR���Ļ&1I��Qo�����ߍ�6�y�����[��B��s��Q_kE��%��Po����L������p/��S+&B���˥D&е���Q2FVFQ�~��x�R[�ۺT�i�\U���STL����%>��?lm$%��U�U/���7���Gԃk��)�ND�9����F��������$�v[�6���K�������oI)�n	�5-gy1d�/�&V�I<}�����@�w:�_�ٖƭ��&�)7h�ŀevGR��/�՚�#	��߷Z��bK�eP�����V[�^���}lzO��T��Kka�w���7/̧xͷ;�Ȕ���,>�N�?zL�?n��4�6*�?�@�/zݔ7�� �D�o����e�\�[�^[*�=+ye�Z*~ew�ʜزA����vB\��-�n�z��YB�xVg����Y5��W=+�2qYr���5�s����u����-�A'��s�vJ�!�\ƍ���%ğ2��͌��{SJ8�q�J��A��+m>�{,6�\��HR����Z�|{�������P���et���G+��s�4 M����{�<i?�PZF����D��Ȳ��A�Lt,*�tUOM��3�co�K�=�a"�ٔ��K��g}��[@�Q�%��W��?zdnN^���f\�х� �¼j�Pـ+cU�u�����D�Y�6�y�ڳ5d�(�*��a�fq_,P����ܼ��t?:���F�sr��}:�6�A�}������DI����%,�����އ6D�ڬW���*�!���=���#���h�W�t��+;:^8��E�ҽ$Mb�����K�j��|x����yKA�6&(S����Ͱ���X��3������*��=�7�,{+T2��s,|��Jt(�*��Z���B�ol}�%nC$O��.�Gg�,� �;?Y�9R^l',��S�"_�e��0�jП@�8en�״l�j �>y�UC]�X^�|�.J����dx6W`}nꊲ5���3�G�ݘǽ��:�A���Ե��^ 2��D��6��������hc��;�:	�����ON�ǋ-X$Dm��ks>�p�����v���!��~��V��`��I��v�\�jj�/�0���{d�o8�ǡ4�ϖ�&'K-Yx�,�Þ_���B�7VY�� ���t���m5]�do`��ï�
K�?'��"���ԓ�G�&j���b�?s%���p��g�?���y��~��]M-�ߓ�O����l��p�mt#���nd��[��°��<���YUǦ��O�ֶpo�u���ݐ�C.���>A��]8[i�_Q������]�J%��"�\y�n��2|�GX�R�G�Ȑ`���<�%﷞+���S辧O��h �0��/�����H�QS2�y*��be�~?ӊ|~�u@]�dhC�0�A�>�G�"�r�Yy�+�[,�Z߹��{_�%I�E8�[�m���E���#�6lvrvL�ƨ�/����\l�f�
���e��Cf�*��},�D���]�;�E�u\�J�G���?�& �d�`��^
��E�p|�27]�U!�O��0*xV����p��<.!���)�P?�6�ѣ���E��	�h P�u�Xm�� �!.Y�f��J�V���Sx!G�N���ʙ�=ə��ȀDz����ե�m?U�N#L�~��K]�^_���
�V�)mı��	|ݛJю�I� k�7��1R6�de7?:�^f�Fp�X�6�	.Mg��<k/�YNM�º�f3�;+�Jt����͌���5��Ɯ��AT��;���'-,`B'*R�Վf��ymW���o�s]9�^��(���0:�J�	�f���Y� ����krr��}�1��iR����k��z
��
SaZ_2�(Q����o�7�r��P�j�'���"؎�ݣ�5���F	����j���W����RL��R#{k�&M�8)��R���ҥ����0zL�{��H4�*VnD�Ho�@"�t���b5�b�9��8�:m�"|��x��e�/�#�@���.���Ah>*w_6�I��8�먣���x�"Db�$us􅞫��ͷ؉߬2�"�^�Ѕv�\T��֕执pXH��`N[|�)���&����D�t+���R�_��/��IvJ9������(^	D����A(��V����q��@�o�n��ɗ��{��p�d� Dm$\A&��\軬��x���0�X���j��
�����5��~R��h�9Z�s�������"���Ӧ�xrӐ�Wl]'Q����|�c�SIN�nTճ�Z/����̇�Ÿ!XhC������'�!xN�{�d����&�/8��yh���l�
����W����2
	,���7�s�J:�Ņ^�O[�'���GHĒ�J��y�u�99��`l1��b�4���`�B~A�s��
���l�H���6N�b��X^м�P.�j�'%����6OE��A>�QAMJu3��=ɶ��;��9�����'�_�ݪ�G�y���7�֋RuC�·�&�K'<��p׉� �z�'馰T�>���PoA��ܪ @�<_4c���\�A�3"���B~8�\�º����^	f������?	2�N��v�"�y��0�?�/�q�4�pɔ�)H��#�mw���[�h�B�ħQ��z�Njg�5���=n>x��Q<�*����p������ۆ���V�Z�N��u3Zg��m�U��4�q�(.�;�_�'0U�z�S��<*C���{뮣�'L�E��
�d��)"�A���b��� ���{��0�*`������3�*-�0�7�c�ː�4�3�elp��g0���b�����Tg��w�8���,�wD�N�mNI1P*O�8QU=�<��j�r�����n��-		�ll�8Կ��'���]�g	X���1[�I�:���̿�I�ͨn��0愍�7.��DwfBVB�Yw�4�W�yi��:�3��o	o�5�p�<���y7���.D�KN�X�Uw�����Ύ,5P���������}����|��Qnw�lvć���f��@Ԇ�1��X��8�&x8;@^�"��雁���ɞt�U�I�Ew}J�F��~��<�{��.�ۏ�N�̈́hɼN�S3���m��5v]���c'�Pv���D�Vq��*_�ޏb�-c�=����j(�����xrDF}�W�1H����� [�y"� �m��0ˇ��]��}�}��	�*^%�~P�Ea7r��T��N�9�{���(L�o\�:]6H-�ќZo���_?�,��׻epI2�.T�r2-�QL�ON��<7�T_��2��>�aȘ�rz��y��R��2�c�n��c<��\��5�Hp�,93��&S��{Y��٥Q#DD�ڤy��J� `��K!Sn�GE��(��D/ ͞_�ӵ��%�G�����A��q[���s]��O��k8g'],C���.����I
�^jD|�~C]�87�?.����n-���&�s�P87�3�DJN>�����ie�k��>��L#0���n~;!.���N����cC�m���(��>r�'���O���(��aʄ�̇ Ĝ�W����1�m�m�b8���z��E��X����􄙃i��3�a��A�AӚ�f�*���K�UC�؝؍�V��C�"PV#�
��n�`n��>F6�rɼt*ԠQ����	�y��g�,��ݗ���q�Tnmݨˌ}��m�~�΄}w}^�r�p�����F�'}l}c͹%<z�����h�d�鱹������ܛ":^��HB� �-�bg�9&փ�5��l�Z0உG�0�j4e��+,
��C\��}�s8�^'d`m�1�6��w�E�$KؓR4 \��	�]��h0R��`%Uߛ'+���b��=����QO>�GZ�,�-"ic����Z�9��N�X��Ԃ�;%��{�ȗ��Ҍ�b@T˿:d�m���C�U'�S���Q�M-�680Ҕ����L��Y�9	�\��?�5\�xF`�Ts���(BLϕEb�Ͻ�}��݅*�v�M��(tF��3�E+�E������)X����/�&�'�
�<	/V��
-+��Y�ľ��WR���?/�l^���c�����O�g~��s\
����̜�Rh�!�y�xo��oÞ6C`r�P~��/Rb��Hl�4��̛�=��-�ea?<V���=��O}k������z)�`0�QtB����c*��n�mI��x�ed
W|��ZVګ����ɵ����v9��?�a:�$�b=������2�����B�F8���w(�"�p@�*��)��&��o?h54K.����/�TF;Z?��f�`]�
.�����Zgt���D�2;��=�T�طg	�j�|�o�N�������� m��g��_j,'~����G���/���X���8��D� ���M��M]z��5&bc˞i�����2P)zX�>���ә��H�ހtSoP���y�Ua����!N֤�_``���&�n�Oo٩�*�> �r>hӌ���Jڜ5�:,�̣�1׊u��n'
��E�:*�n�w��ޠ{!�Z0[֗��>�i]n&�y���ͻe�<��AX�0d������éI"j���4܁���{����S2�_P� �E��\R�(;�P�iD�p�6?�v�����9B��Z	�D��M+kuF����6�%@���N�ReT-V������K�l�k��o��Qr�#
L���= �o.�6�.��*BeU�|��_�`��+��d�㾿�Y�������l$����V�ˣ�*�jiA�V���1�v�xG�y֏��-<Rf���ҿ^�Ģ��B��K�߷��QPy�M���BA��M��׏c��393���U��Ζ:`�����9q��g���:ۑ�ݨ���?���:�TN�,�5d<�Ǳݚu�6Ɏ�C.��5��u�˙kl˴�%^qk-�"�L�/�=���h2�\�iT��<��j��$��6�3:���"���@��_�m"����n,�
�Ƌ�#��9;��/�KN���z7#���Ĕ�o1de�vPt��[��=$����"Ԉq�	�u���޴���L���ZWl^㭼T��6R5��2HNH��`�j
1˙�{y��v3�I�c��x�۹$1O�;��?{����q��O=]V���g�M��|�f��[#I5c e�e�zDA�����g���?��so�f��
ە-�k�O���!XԔ�ЏRr�I�i`�r��?�Z�u�J�7�_�������$ �
cI�Z�+�ǋ�+ٚ�x��ؽ~/�?���`B*,/��z�Q5��S;��v@���kЄ�	�&u���c��am�ֳ����nTd P��1DmplNf�ZF�W�:$q�Y� D�L�5�y	�.�|�Ϻ��H询���j�|���m��[�'��0��d銲�2����ho� �C$V��[1�G�n�MO�l殘�F��<���S6p��hbo�o��z�/3����ȝ�.~jg=o��.NŊ��_�������A���K�N�#r��*� 6�1!h���	���,Q�K�~:�K��ռ��V��;D������s�ǜ So�j���'��H��Z-浍�����<�yK�=����ܮ��}�M̖��$t��E=Z�z"|��>Q�p&���D*���&��>]�%rP
u���R[^���;��UKb���} N�{y���7������hQ���d`C<$�H�0V+d<'T�e_mI��g[o���B ��G-B��;$2��!2o$��gV�;6K��b������-s:����}L��.R�-*��T����Kr�h�5z���0[�@�j)󶒢D�(?���>�g}��	�V���L<@z������!� �!_�R(K��<S�6��@Qqa��`� ��8�� ��U��N�I6�d�M���]�tn�C�ᒝ�v؟Lc@�n½Y���E��'g����I兖�h��6VB��v�Weg���ٺ�j��W{��kz�q��Y��N�XR�U~������H*Ve0� ҭH�t�#^]s����?yy��q�R���{�!�৏!�C�b�6��׺=D�Hs�dj�e%� ��+��!h�s�vr�k/9x(������+�0�L�H����]��̍�C){Q%4a:,����d�� Հ�XI�D�N2���,v�/],�ư��:�d�a�R�Ezg�'�A<��T&�'~E��aB{袿*��"� H�����5����3��$�yn�i(|��B�3�'�|�͆��s�!�]D\j^H��dD�~:#�����
���� �:�."[G�u�4\�#8J*ش��WC�j�ǐ���w�! �FH��N���K��o骃@.}J���e��&Q�����-��ҙ��5��^W?N^lg�S�k��@��F�_#\�76_e1Y�1���Me�}A�5v��4��RӦ?��4�d��laBs^}P��D�[@.����7�\���^Q�� <�6�I5T.*��� �pT�p����buJ!%?�#��|���l�=Ј�M�BX\����TTYY���+hp��o�Hf�kf����:H^�.�⒎LR�zs�.B��r��s�2�-!��(W�?g�.;��N��91_|K��F�o]؆�A6��I�޾'��`�Ҕ.W�# 3�5�l����p�_��kϭds_��L@ea���~�����ď� �E�u�5��2���Q�Ƀv��u�ʱ�4��2��)e���YC_��?[�i$[7��T0�%v"{cڜ�a8��(�gϷF1��dK߳{)�ȋi���y��dA���8��1^
Ai���*����9w��i?��:V���HҠ�s���	��у�ig��d`�ɕ�C*v%��uE�`#w��N����Q��a�U��Ҿ��Ŗ&^%~ l�S�t�!�E�O�q�@�Z&�E.�Z隇d_N��K2����j!T��V$��rʌ*��5�;�����JX�������ՂN�����ϗWut�4�-����d��oz�-^J�{��NA�챺�EP5KQ�bH�˹6�������0�EJ��a0�^�����&��7R�;��[!ES���W sVF|ۆG���J�@��
%x\��c�(�[�]"Ԗ$D=�$���d����E���1����))3U��X��t!emޠ����_b�jB��
%?�槌��Ka�p���>��O�Gi��߄	�q^9*�d����-��Q��@�U`d���/����S�����gs��p �V���4g�MSu�vIY=l|���2�
j��
����D�{M����"�D&H���5�	4:d;.���~���.�-h��*o��ӳ'h�|p��$x��3��"AR~�B�o�~1J���^
0X���|�x��eԎx��,���Ő��X^�{�I�Sji��M�P��]�e���O9ß?�k<>۹u��}�u8�̃�&]�Ҩ�=��v3�7�P���k��B�wk�}����_��0�_�n"�D����j�aQV�/��d�*�2��Q=.)��`��?F�[�jڭ�X�O�-�x�E����ȓ��Ŋ,��W�R l�����5�~Q*�W(��D�,D�8��X|�b�P�k{G�zpB?���o�~ė����E.���J=�5%-/�U�]5��q�A����6|��#|"���x�3e5+��{��.wZ���/��*X�������=��� }:꫓���n�y�Ӑ�*�@u��p C2����1�ؒ��&�BG��򯡀�~M�wSu]�qI��M�+��M{i+��4�)^�z�A0�Uh�ٞ���
��|wi�^�L"����@2� ����wŧ�Β���/P��)^�t42�c��?n�[��ͭ��D\f�;������i�v\�]6�|-p�'�;|���(mt�10�6'u��k���M��݄�U�3���cD)܋0�"�$�<ۼVN,���G���@�`�$�c�`��`�벋��&��b8`zN��1�N$���*�]���.9vi�ٔD;c������g	$ݟ��V�:�X��[�q!X�����}cݻ�p;���s�N2!��߽��,�#*1]�F�l� �9PĽ���k^�j����,�>i�$��v���銭�qH��L���'
�����Bu&9*ڐ��;�{h,U"\{��_��*=�'Ǆ���:+��+�/����[��M�4+)	z�3�I�A���,_g1)�@o��_�p�;�#-�&X�n�!^���� 9��b 6.�0�����L�:$uj��0��:�l,�/����z(��/e�A���5@��ޚ��)X��X����U�C�;Hģ�f+�]�
$\���� �t�	8$
���s�v�S&?�[9�>�+#���%����/�ػ<��!��K�3$�2
>���<S~ �L�"�9�P���9H����5�_�L��
#q��N<���}xs�B��2�?��0CD�8[M��vO�䘌 ���q���iLa1��~�Fu[O���z�^*��)�uA�7��{uC�L�l)��a5��6����!�'���&��l�n���K��Q�i�g/�/�H�5��6��}�ٶ��朰�:n�pj�E /-�OtB̸����K�뤂��KP�1-�1sr�O=��<��էP�9�93�±ޛ��c/TfNI�D�K��m��6,�/��ϡ�-����ׄ�B$���s�؄\��s����g��5�.���^��qH:�˒�.4�,Zz�F=�~�Ԑ;J�H�N��p�`-��w�k-�5L�H�m�@�E[��`#-����C�G5maߘ��� �@ i_o��`?�����a�u���g:ԵC���v�ӬI2��������;9ڋ{��4*���(�6hgw�����C~S����y�yK�WTbӊ�E�\��p�Cۍ���<6��Sa�Bv�-<%�q���3Hf�tq$q6��̦�����c��$�\�P�=�Y�쬥��κ��yǋ�韥�l����4�8]<���/n�f=u��E��Ӳs��������+A��[>ޒ�/�LѮ9�O��;g*�*���V���k� �шx*$�_S|0�|8�࿊'4�gDŅ8Rl��'C���	a#�ɜ&���g�i> �ɫ'�d:#S-8V�����I�.��֙�|eZ��>
,=����hĕڧ����^rL�
�wH#gd��ЯI7J�m[�Ԅ�|����8֗��̚�\����WÌ�;p�؉��m'g��V�\D�,.�X��s��¤1�^1�O�}#�|�Ŧ��֋�� ��Ƴ���s��r*Yc��~��oPv�ib����ۡu���0���5Z��*2�ucb�Kmft0��	���e�G��|^���UÐ%q���]���E-q`G�W��]�l��iH��®�g~�eL
�p�K��j�.pr'Y t ���g�=���Q+�Rw}֜O2�|�U�������>�?����o^��b)̷�3<�E���R��96���U�#�H�X�h��X��Qq�ٻ弸~�5ƪ����T���{,[���BM{��ǌE��.��Mb5��$�}���ٶ�obS���!�r�=���SI�(}C.!�S�9`|ٴ�~�4�t8�¤_($���6��6Ƙ<�Ҋ�R��@��N�=�	�Ԓu�"��i��S����y55/`T$UՒ��8�2�C�#��;���L�5h�V�a����C9���NZl�_��.��a�C��+,���#[�r��X,�8?�OԊ%ELpc�!Ckqy������8,�w;H�������:k�F ��wv��.\��w�*� ���sr�Aa�lмY�w�����98?������АB&aR�0�U#��\�cN��_�u��瘭�����}�����g_���5�D�2ab�������y�.Z���>7��Ed't	��蝋8�+�	�Q��6�f?�+�Yr>�C�|%C�2�j%�����YD�^�T�N�P�5=��v1���+�sN���V
#u ���g�N�İh�i��� m���sd�K�%	�e���w�z������_����)_X�_j������yܡ7$pb�b�ϣA�j��U�%�������OFFhp�s�`d3^�= ����Ky���m�%�z����^�_86x��`��7T.�S��Q����#���^gS�ri�Т�ID�uR�xآ��')���΁p2-����T<����,��߁�[�����l4�+���