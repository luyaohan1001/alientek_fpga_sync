��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���������1.Ձ��/��٩�w�X��`�eJ0 �	�]���>���9�G��}���%���˲#SJ�*r����Z�)@����x�P)��i�6���1��Ϥ��9���V�U�Xѻ����Ҍ
诀��
R-�>_ǳ3�>��
	��Ŝ�����P����p�����̱u�ѐ0M��%���e&#JF�sCQ�҉���{�[�I���g=��!�~��\�?�^�R%�g��e����1u��ܹO��&��)s��?�.��H�!���+�����l��~�sw��t�SؐYPJ��i<lw��"W}�t� S���0��p��Dէ]��T�g 8�Z~���/�1���r�L�̩��J���l=#���h���V�}���C>s{\��9n�yG?Fn�C6�T��닧B�/,S��f��#��>h{רػ��3���%K7R��^�׾�m��t�4\;�ja�{�}.|��:��+jh��\)o���D|�<>o6w:�O�����dr'���A��B%`y����a��w>�7�����w�q}ZП���B�$o��2������{�EH��N�#nԇ�dQ�'@�6ت���n���U������5Z�(��[.��I�+�n|�Sl�E<��).������95)򩏶070�a�X	@f�<X"��W=��L�l䫫+�A�A���-�3����KA�7)��:�>7��P��*�Lٟ�����y4�T@����Av@�-�\35;�.\��G���57]ά�;lg�	��-���p�g!�d��l��❯�,�Cwx��hx8b�.U*��CQ���57"���~ۧ�A�w&��ϒ��ce<h�鷳�#<A�E����"K\#�� R^�з #w`�j_O�;J�8L�������	�;y%���t~l�4Eů���Ti(���
v`�Td�y���`����,�b���zl�bb�N� `�d}� �yY̼�Z���XCꄶ�}4�8d�瀲��Y�����q��j���}�9��ǯ5�ާ�	�żN��x���~{��FKX�J(���FLx�B�|XNBD�bf���h ؽTƴ��z� �lG-E6)^��a3�N�3q�n	Eu]Uﮖ,����>��$�ws-��QvC�t��I
(bӲ�yY󯸢haM����X���R:�W�#��;��@y�W�zh%n�L$;����[`�3�;R_��$E�����^*ؼ�����^����'ަ O~D��5o3��Aj�m���+�$�a��O�A� ����-B�v��̹96c���7$� ��r��)u:p9$���B&鶰��)�2�:���~��|�Ì�Y���z�i1)>���8�,��n�W���8���$���Ʋ������j���Ry[���߭�&\��^e _��Y]Ѐ��ӧ�߉CO37>��|])��VS���+Ҩ��unw-q�%���Vsᦍ��d�n4ve����M��q�!�>㞦 �ˀ���7s�Te��0	�p���2�yp����u�w	yЍ�X�g��/h��i���j$0Մ'3tts%*�H�������M��GX_��fs]���8�ޝN�X����ѽ�-��X,=+���1w~�Z�P���:��|r,��K���"e�t�G�^�Zb�E�1��J�/F,�FG0�R_mk!9��W�K�So�&ʩ'��p̃S�	"� ��ɭ�����x�
׶TQ*��s��w��ɷOZhjE�y���[C�K�V&'�	�{Q�!z�ȇ���%�!X&4L>aJt�R6�h#��<�[}O�2��w{�ʩ��5Ԣy.����b&Y�koq�?ς�A`g�l�Z�>)��2wf�LN3�]�ElK�9�r~���)<8�(�u�R}�t�I������8iv|�c�&[=�뻆̓ݠ�ӣy���Y��\&����`80
"f��B���N�*M�E�3s�B�t��ĉ��ˌ{VA��,�JA���fl����d������PgC��V��K�d!��G��i�#�e�m��3�鋡���ש{C��rL�l����[�k=�y=�������1�3;�1�#H��(��B@��D��0g�[�YQ#I��u~��U֐o[ނ%c��d��{�w7N=��t�p`~	���o�a�ūO� Ӻ?}�5��Bdh��+��s4q��^���տ�|�Z'�/s�_j��3Ӟ��A��C���4g�n���q�_X�w�[�|7���pӋw�yrT�K�A�EY���lpq�|��_�!��������[šTD��5�q2�[M{���������3�<���5Ʈ:�G���m��Sr?"/�J@��M{c������KŃ'�+�T'���q�rXD?�>�_�I5�,���ߟ3�f|	���H'�b1,��L���BN!��R�j]O&�W%(��4ʜR���/��W[�.uY;��F�\�s�M"XO6N7KZ	���qM�18Ԁ*%�&�R�z�ܷ�����)��f-�Y9y�$�1��p�w�_��DKg1qZ�]<m����Ҭ��ܚ�9퀯Y}D�K���ܨ�M��~>/�6�* kn�n)v՛0�_&1N.�5׮����)d��A@M�����'0ER��ܕ�n�6�ե���Nn��~��7uI�v�'���]��"!�Hqv�v�1�����
�._�U����M�(���X��)'��H�*����|L�� ������.�cK_p���+	1Z��%��8r�`���;G�n��2[�@��߸�{��nI��m�������3g���M�	��'��>�*U��`a5�m�7���	�j;:e�z^:��:?��'�L���~�p�, ��5i�Q�#�LG1>8��8�o%Jj�T�,Ю 5���Է�f�L*��k6m��^;����߾�߄YҦt�O�a��ƹ	�$n\j�u��.��	�AH�n�d��N����"��TI0�΁w��#D��&�W0˟Zi��w��%�h�s2҈
�ЉP2����x��{���&�8���.�}��BF���#��G���
��i�W�������0x��t|%��3��_�U�� �q?PK�w~�п�{|ML��@��׿ݑ%35J	3�ǁo��V�XJJ~ ��'f JI����Ȑc�M4�aaVº,�D7��;Fd�'fJ��$�]�Οf`KǊ��L'9�]_��.�~[�C����֓�M�σ�+�j@_��7���ӂ��EjaΣ�f��|O��&ngU��A:o �s�������2�q;�1�"X�����3�U���]g����|�d(��=����k7wr���B�-\]Y��w�'�&hu�}6�*��m���[m�klz&�cDD�l��|篷���'&#����$h~9�6p�4���6q�qU�AtS
�2O��S��s�Q�i曜�w���zwtW�	ܼ��90��{$2Gn;�7��ݩ�@����Ŝ`S?R틊�R�@3d�u5�>��N����o{�_fNYʡi+�놡�������x���R���TJ3�5�S�)�z��g%�G%2�����ҺNP�����2��܊��B���z y�m���J���,�䞕'o��a�O��Z�5������ x�4�K�5S���hG�>�I�,��"�Et��ң�;N3������a���tw��C�3�kUv2?ɲ	��f3	.��{���Zt�B����p�+��¦�<u���OБx�b����vt^QA�;���%׫���-a?�m�m7�h���]zd7���E�O�hǙq���l`k��[h!Ćy��� *��0��\�K��(�ב4luǃ�٦��lI�Bў�4�u��v�E&x���EU�9��_��~�D�\�Ie���*�h�����Q��l��i��`U�1�Z��O���Gx��2k%��,��A!s���ދ�k�j���RG���Kno�쑞��雩OvDXq��X�3(!bq�H�+zqqnO��l�/�#����q�ќTWTJKT���/�/��;����@?�N��:��i������6/�p�kd~G���_fC�Fm�����c�/��6�>��[�p���pn8C��N��I��?��P/��X
�w]*�)��?��gE߲k�Jۼ��P8��~Y�C�/�r'�� >����X8G��m�m��`�=�cb��I�_�Mp�����8F�޶�P5(%2{����)�SL��L&V�K��T�Kl�Hiz��T?�f5鹙��0��s��CЕ��a�޵��2N� �uR���l���~��2;�9�`��x�s���#q�3�%�2�?�����������L��,9����s�5��D7��3��x����ˢ���fwo� T#��'G�����Q*I"��fZ5�u��q�u��*!ͩ�$˕Cd���٠���S�O���R1�`�!9���Gi�E���p�����53!����nv�b��j������*C�Ǣ��Pg��:�_����I@W҉���H��*3f�����/�!�-���iTuN
�`,��F�Wu��)�E��5�LL��|�2�۝�C1�� �-��$��\/����pn��-Cg�i��Ƥ'��I�YT����~E��C�n�F j��0KF�g�����Y�(�em�B�!�%��ƣ9b�nY̿���ʤ�uy�;������{���R�<gaz�T��Q`�u����I��nY�.��s�ΐa��+���Ll<6��bI�ɷ�4Զ�,n>��}N��oE��
|�!l�Dz�
LV��$��vl2Jn<�h1q}�im�wЖy��%�JP���L��3��/�E�s�c<�ٚ 3UM���ͪ��J`D�.a�g��;�Rp]"��?����z\�Їa�5��=>�lS��R�v��$A[�;���qǎ���`��H��,��K(t\�"E��_·�Ae.u�,�6+C��PߝYt��1�H}�R �dtI��)��t�smE&T�ci��yiUȦ�T4��t�3�a��i�\�� �_��¸�Ʈ	Z�A�8�˻�0G�&�2�Hd��i�َR{E5#�wWH'-����&��P���S�;TO��X��hE�T
z�}�J�?G)`f��9\e����q��C����k�������X����C�Su ���a�i(����e�&Q��k'��9w	�q�?�ytW;Ō㉮��W����o�JYXSH�J5D�6�����@�v�j-�~�*rV�<�_[�1N_t�=�Y�ܤ�� s��Y�c� "�e��Кa�������l�ec�O��g"��zn���Y���g.:�@�`e�L���˭�ێK�k����Y9��.*�ɢ����uPi�k؅)V��<�B��I��&�G�]�=�l�.籺"4}@D���s��)��e���&�i��؃PRV��Z88�N�"%��WR�0�a�u7\X*~���1?:c��D�]��J e��_��K��E @�Rv+Q���+��"�V��.?_�&{�ޯ>TV=��!�%<R8Wы**�;�?_
�Z�k_~�;	�<Oq��~E(dN�Ձ«Z���8��̵�G���b]�TMD��;v.'�c�Ô�_�P�ld�A���z<8��VA�uG�(���S�7�]���Е[T���]fԯ9@��ڍ�L*����Ұ�����>f�������<��v,J���`�$o��(�%	_��)	��5G~gTru�Qmq�(�K	�W'�_��35���\�w����k�;n$��0�gR&�d�m��&�����	��E1~�h4D��{���	2��wӿ�,��U^j����?�`�*w�O�⑔A���^���HK�N�V$�	�f׀�_�NK}:������,��`��/�6��-Sɷ̮Sv����J��e�3�I5����t^��pcѺ�a+�+8h{My�K���ž{�Q@~M؉_��m:�`C�t�sx��h�lg���2�-���(����<��u/Om1F��u�:�WGb�bc��	p����V>ٌu"w��Q��ѣ�̞\�8f�n��� �2�35f��P[P
�_� ��K"��X5ǂ�b �隄�ցZ���M�-_V��`A4
�sd�y?]���)�{1���g�+M����Aa�#ܼޥ��v-�� I�S���A�ޮ�Q�X��2йƕ�c��c�$��Γ倵k@'����'���W%
��84\,�$bp�2o�\�N9��N�\�c���V��5�����v�����E1����ڕC~��a`�SP�Ց�Kw��	��l6UM�t����SH���g��-�GT�/�8�r���2�T7�rS�n�kƯ8���$�J��&]L�����줾�F���6�M��	��Շ��ld���b�6�b��xQ��o�S�l΃��[ae!�u(�����1�3نcQ+B@�����Vk\�����! ���4ʽWd?^N��3)}�Q�ͬ� ��+RIX��`��_&r����36��L���.����}��f������CY.c=��,Nhf~Z��ˊ������6}�SE�Q�>�ө���&����ê�rڼ�zu��v�y᧦�^s�x�~|�]��H8�}`c��e򢇏YD�A3v��f�o�%��L�v�UN���Qj�Nj���2R
_M\�Lc�����ׁ�auӎ����c0�[*���n����=K#�~5tuv�k�1�
5%�.g8"׷�<9�p��ћ8�AP_�kV����,=��S���,Zh�uW�WmW�ȸo�3�"�e̓��>=�Ye}	��!�@H��/�/���VoLz`-{7�e�@����mmT��L��<��A�2�a�u��}΋����E��\ ����1~�?��d	�o�k��*��l��A�(#��e�'1Q&��յ��q��a-�!��Ԃ�?�W�vdbC�uw�V������F�4�D�\mp���^Qm�!Ym����W��y�۱���J2z%)Rg�n��?~�a�����i�ݯ�Ac�@�_��V��}�Ve�
>�xz���|=>��0��9史�����{*l�yp\�/�8x��y�;�R�[���z�s+��R�ԕ�bV�'�9g���;��h���i��/�F�ĳ�8UÜY�^�j	�k?Xs�E����
����b�;?�e��+��J�Cc�o&"+>�(U(�i�M���f�sn
�3?q4Nj`j��rE�qȭ������J;'�]��V9o�q�!Iz��7Bz�{Ahd��$����T�?BfQ�Sp�9˻�#$U�!��1�3�ه�&��2P���Vw90 x��y�M( }zBAP�a���7x�$&�5����d��wA�c�HI������ҏ=�s;F&I��Es&�w�q�7��R��r�?�t�!��xhP2� F��]���n5�OAs���n[�[�ԅ�:��FpCm�a9|-�T*[��2$
��h#N6[_+��5�aQ�V��_	�g�f ��D�K�Ix�I������T(���s.|�u���}�V9�Wj�Ҿ�I.�	E�"�t�	 QW\RC�B�9�a~��yt�W�����p �:� ʯI�_-��.Z�I�㔆�#�>��� �n�caWj�ct@� w�߭Z;���2�&�T���s���ݺ�J�e,#�,����9���/?��2	mz/��A�bv���f���;�'�'c��k[+��Y"�ӓ���T�@?q���AX���-	f���Ʀ�-�_A7�%���T~�����`y�R71ʖp�X�yD���K�����O�O�����h���p,B��
��Ȏ3�P�����i�����S'��/�lL�
�e�7�5�d�����P��ЄBn�X28s�0;�8=�=�Z�ݝ��d�U�y�Ǹ�-!]G�t 4y����9��-��~�EO��x�	3������OӪ�8�k\��#a���o��6��X6}�	6���n:�qnGQH��T����F|�t�7Ђ\�=u_e�O"B��h/����R������؎�W�ָ��P��q�Yy��-A0�,����Ⱦp��8��F�ZY���ș����n��	�������t�n-w��̅��#����*xj��#�Q�M�'��%��=q����>.בP��VF�����12ק���H�+��WK�o�J�kI�%Ri�"������{®[�0K+�y�}�1��`\�L����䊫a'r�tX]�O�8:�ϳb�|��x�5�'�i�w�N���A�Z��r�0&�I��Apt�V|�F��B��-0{M��LT%?�G�zJY`�|$��Ah��P�R�mr�ayLr��ݱ�k%�b�K�7K�z"&TΥ�ۃ�#�I� �ST�Q%ٖ��?�z�[b�tW��Ɠ~��]]���I&zq���S���D��u�&��|�ޘ7�ؚ`2�#�W�wc�g���+��4�]g�x!'Wb2\w���I��]\/����^j��Ƕ��cm��� ���;�z��D/�к���O�������,�d�g�B���Ì�ss�}ۘ����z$���^br�s��1icO5E����<��^�/[�&<+����|�s"爪6% �?u{ML@nn�zZ����,�
X�8�UBx?��F����S���#�81m����Զ-Oiv {>,Mp�;�߄��M��7VJ��4����/���{v�X�|b[Q���0_)�_X��&��=��H!ڴ`f����X�H�C+ �����nx�XW�Q3�O�s�b�G��nv�)�s����9�Y ^����FL�<b���JrW�s�x;a���������}e�0j�Mԉ�C�@�p><�a[�e�
G��r��-{Ms��|H�����=w�by�	����I�n��]�<�LWO�2$�j?)&����)ɼ@���5�ug�eu�8R�q���B�K�ۡ(�ǐG���8[�Ty3�{�����dJ�Eb�13ؐi�Lv:���+;�������fү��e\V֠vW 7��)heF^�+�����=x0�����X="Z�#�6��x�ʪ���am-�{s����E�Bؠ��u��j� p:�	���jX�e�%xQD�+���{���u�ޤ���[pU'=x�
>�d���e�&�)k�&���_60�,.+�����eD.�>�!�K5Yc�����
֠?�����W��l7j��Z;F�����*�i�&���Zi��yy�uvI�W5���Au���;HlEg7hrZ<�yj���(�38֥��n�DM���O��C��*� ����މ<�*����iZ�v%!�����/�;���ӯLe��bT�T���`^���Q5m�h�4��~��F�l�W��rC�����w��Xr�=�x��N�J,���5�꬈X�RU���|�~!������"��`!���
�I9%"=����b0������Ќ�m'쓲��wi$�������@3�o���$��vG�ܛ�l�!7ƶI�!�+�o�մpȄ�<|�]M2Z8=\f)��I}�x�إ�W����v6�m�@����w��'�=�[�r1�
d1���Q �U;Pǻ��)'�눵j�%!�K)��=��m�o�n�2�CBH��V�>~Q�Plsk�R�`�h dC߉v�2�f�;��<�N�ZʑqVޅ1��+a�j�Sw��[�rr8F\��P�N�.@�����h^B7P�������3�tG8Zh�w���sJjeXu���̾�5���mWz@-�Р��f?�m�$F��Nx8O��ċ�^��r�%$2�9�zJ��Լ0s�4`� H�5m�p��	����O.�FI�eu�y�č�ʆ��ЋȽ3��oh:���{�n�4[)PgZ<�.�c��ݱ��L�(I�ۮ��ƝZ�|9&�.��-O��R�4wV�'f�m�m�LM%������N���P��xS��/�=�0�G��a�j��+&��u���H�ݘWc�"�t�%��w��2�+����j�B͹��i(	�ҧmS�蘽QD������bж�?h]IC(H�$�I�t������x��9��.0��tg>�c�X)}�$=�xh:��E;�=9:���r��I]1��Y��}i�P���P��(���n)��ǎѨ�0������4a��>�{r?Es��w�~Ln,���V�_�*�9u��X�.�7���bT7g���C�S����I����O((m��h^8d�[S�Sk.����OL��T�9�l�f���]�!^m��=������+�?48c�`��+�eu#�x�!(�a�.� v���4����$�4B}�+%�F�erF�Uގ������qK�(sN<�p��JW��>��9	��Re�TU� 8��2�t�I[Lc�?�݆"����=Ŏ޵��-go.*s"X΢�H�/����|nN�=}'d��(�]���WM ]���"�83ӛw�8c���=؉g<f��NK&ݝ�b���섭|`b���N������D��;A�ٝm>�ĘT��£����< z�Յ�@��L��L�Rd|6���Ӑ����J:Ǆ��G����J5-J)��?V1���y����P	B'C��R�����oda��E��"R�WD�E$ϥ��9�~�����#ʴ1i�R��MV���e�T�"Kv�c��j�9���'1��T�y]oG,������y�m!����ƚN�r�3
��*?�M��'"��}�j�6]�+�BkB�o�kA��d/GQ@ۊ0H��(+���S&�|�Z��g�G�_��w�j��	��UHh����R΅,�_��ܨ�%g����9xc�w�3�/�}�(�ԏ� oݶ�\��t���̴��)Iү��{U��'~A^�n��.Z�;�ǚ�Q��dS{,�� �N[O����<E-m���q�ekB`0e��{Zb��|�"P���%��!@�m�V.l�7�	�%�!?K4��@Z�0Z9��x�r�>�<"�~H�ȸ�A�#�zI!ElC��kZ\Y~�GF��Y��]M���qf�L��}y�w�@��ی�����
ꅶ��C��Ŧ��þ��.Vw�Sb&�ϱ�IX��*�q�K�Q�-����,���;�^��=�>u��I��xF8³�����R�~�O�2C��#6�޿�̤\��߶n�9`�<�do[��sS�)-���Ј�U�#L$�}��N�_���GŁ����S(p�W�MGPG��v78=� ����F��oK�[�@l�?ɠ_$�u6�̘ʿ��4�8�.���>��ڭ��p����7��/�q���Q�{�q��
\|�<��1ٓd�_���컋��@�$��yѮf!x�^�HT�*2M �z��V
�����t��ß��hnX�6��!�7���Ni
ʴ��h��PVo��򭄘ǩ̎HRp���@_���������A���~��;�T�2���Țd��t�1��e�D���H�s"��	\�i��x�^2�m[�m�_�[���D��u ��3^\k�cj��#њ���@���/P��2��i�U8q��ǤK��D�n{�RX��!s���wc^�OZ_W�%�����v �TU�K^�DF�N~,��&��YQ`�ǗV1���;�3D@���a@L���tO̻}4'��䷷ӎR3jޤ�G\����������D�m�O���� h��ȶf��>��<wpȏ�2(�ַ��^ �b���ne�p�o%j�
U_���s�z�Vnw�"پ���hc��1UyI�DJ@�T��g"��F�l�2��
��0��<���%�Ɛ)C����.A+Q:F%�0�úJ-��kb���2�(�\�"Z��3�RNaÎQ�}�!
�A�"�|��MB�"p��VN�H'�p����Ĉs�	u@�T��4�ߠS���b���:�@)�ۘ4�D��x���v[�����e�Om�����X����s�B0���Y�7�]rq~l��?�@y��:8g��B�n1�关�l�MiP��>��&�����,1F��f;�e��z��nPh���8�;f����'!ô��,W��4Q,:ɜ���
���1l~�z �Q��]O�=����	�f%K'-��!Ʒ�U2l����n����`�qB>�cj B�Ly�����@���+o��p�o��&9��$�&9�F3�+!�~I��gy��r���"(�����IOT�pR}�̚ܢG�G�(�;���G�w<ч�S�i��s��u��� ��:��������QCӦ����;�3b3H�&��ٞ�*� �Y� Z�nC6���a��.��9���O+�y�3!��^E��ݸ�Ȏ�L�L�l���������貽B���q9B�C:j(�Gd�h�����\���'+sR���7�["�L;�+�Z6�dѽ�Ú;3�R���]����^�`0��;p���TZ��l�f!n�ُ����,P�p��顄u�Z� �e��:NQ���:�K��F.��BHt;�	�������+T�_ծ91�HF8_���>x,`��vɦ�m2Gk�D^�|D3�w��zो�(
X{����)��b:4�>Ù�e6%Hw�W2l���������k�;ND������d�(���0:{�h�$�ÏZ������Nk]z����)��7�a�v��6	r���]@9�~���1������d��@�جs�A��c���w�1��B�mc(���R`�H��>JJ��>� �C�@����T�6�.o�]a7�����T�G=ش�E�G�N2�d��|�Aٴ�E{tJ9a�Y�©@i~����Q�X�(:`a5\/j�G�1�Q�?ah+���{q�HR�� F��d�֏4�a���1��(�QS'�%u��$������0���"������N�7&X��=Ňw��z�;��"j�k����dF��r`�yu#��ٞ��gL���X�@3�Ѱ|=i1΍ŐV�:�cm�F5��:�]�?��۽�b�!-Ï����tC�?V�GUm�s^�߆\*.ş�Y
�������2�	-q�?i��cW+����O�����`�������#Á�X5��ǌ� P(q�%M1�D��%��'_�N&Xm.5��fkK�9==���<�(��W��0~W뙘�#P��O�T���ϊ�*�tP��_����)э9?>كG*��~7�!9U�=���s��_hCJ��!ƿ�+��6=���2�e�ki燡������-�MlE(�����q����:�0|� _���i��Nہ��O;��v���Ń��b�I7f�Pf��X���|�!qu�t�%��A������쾖㦪>�_�!#�&QG��\E�U��K?Υ��HgH�b�A�y[F�Y`-�w�Lޙ_WH+I�_��0�s)ʔd�����-`U��y�	��vk�񇚱:ӝL�Y<q�%��W�M�sך�p� �A�g����w�ڡ3>��*q�uV��9�L:U'��)�W��ufO�&;ґf's�����ex޴,z��>���'0"����u��iSK��Tj���$g�ܗ�F�p�t�Aڨ�8����1Xă�;.���/�3��p��wz�%�+;S�y4J��ש�]_�(:�&����>��m(�Ø�P�\)6&G��q��Ҟ{|ǌ�ܿ+�Ώ	(�'Cn1cpw�(�P��􀐳רZ�y;��:h�D�D�Ya+�N�i�5x�9'��X�e�.����u�k��z����_[�%L�@}J�.N����ʒ��`st|�#�A�9�0�U1�d��W#1/X����%iC��%���Xy�^�%�jt0�}���`���Nӕ�э��Ƿ���u�)qƦ��OE���m�j�����m���;����]Kb�m]a'�Tցv&�Qe�>�k����������J�S�S14C���1���ce�,�2	K�%m�!1O�É/�*�	�`��{CTf,�"�� ��s8]�a�قB?2,l.a�|������
��DG�R����ӑA�Ag���;�Ԓ�k�L�H�K�'.�K)g�������Ͷ�ߩ��u8�R�|ߔ���)(���<$�q�CN���'jc0�$��Z���azFV}�7�$S	�����K
s�K���8!nw�q�E�g�����/E��.C��se�}��.��Z�n�λP-�; >�H�����O;�t�����# ��X��r˫�l��}��݈"� h�(h��r?T�������w<J���ɼ~��r�r�%���
�2����[:Z3t�����f���m�
��-Pϟ^�5u:�@�/�BH��	ݽ�	���x!�Rz��]X^]�Z���T>��(�)&
)'�X �s��3rڋK���t�)T=II5�q�y5�H��w��|�=�}�U�^�)ĿV9�>#,�����<w3�A�Ԫʵ��,��J��i���;�~fV�N�DI--ϼ�0S�쨷���EoL�o{�e��&�,1��[��is�J]��ֺ��O$MF�O;=7�jp<�f��Z�y���b6.	p��Y7a�d-��/w�5Q>� �ۯ�L��iK��=픶�l?U`C�Bȍ����[A0�
!�>w��N�G�=hc���2]5k̩��-{Ъ	/Tp g����W�3�S]Z.2�Kbc�1&gh�<<��%��ہ�o�<�JY+���&Bv�аc�zWqaN���^��[�Rn"�ٌ7���M�:�4�)���0�}4v|��̠�ڸPL^m��t�߼���� nH���E*��{�~���ʜ@71z~�DJ�(E"��nI}m<�5�/�~�!>=�|��f�ш4|}���"�7"w�����.B�$�\�7s��s������'�[��}��k�S�Q^O6�)����)���5��}��}�=��~{�;'�}|>�h{��׭�;+������SbMp��Pˮ3i�d�P��!��m��bhzv����{�Y3y�~b�v���
A����'�-O�oXX�_����p{��Ӭ�u�C0E>�eo�P���Y��Z��޶���B��g@�������/$��}�
�.X���d@Yg��%��]f�T��6%�� 8@u����g�@ӻ/��s�d@j(i�up\���A��{-��p|�sj��Z��by�_w{�^Rq���O���y��H#����Vj|́/7��[Q�6��	<��c5sB7���D�S�X�SNA$q�ٝ���/d�Ex[�V�gqr���3�"$6P�[ xL7-tq�xb�����MT#�%��/��Of��Y=.���-�4��Q�b����gFVD�q��>��^�p�[�/�)������ٳS7f�a����+�-��)�@1�x�����䬭�Ǭ�	�S�'�� �Qxj��	���]F��v��e�7C�(o���ϗ����Z]ˏ�>hsZU�����3�����=����h�>�"��<c]���Qٯ��R�,�l�/}�`d����;v�ɀͶsO�UʕN�j$�M�?�p�HXwA���
�[���g���>��K��{
�UE�p�hot�!����ԡ�4Y�H��]�ŃϘy�0e� �3r���1��H
k�;���Ez�Ź�ç�'.���bG1�J=�m��yI�m��V�β�9'p��?U�I"ұf��\�q�6^�z��7�P�+��h�^T���e�����hp�*��kD�%+���F�,�h�@1�(�w��>�� ��ئ\Q~M�u�1I��9P���C}p䤋u1�X�7ʹ�\�t��S�]�0��ޚi4�C�#���)G��I�l�=�A��n�\���C��T��r��V /�*�J�Ka�B�O#6�?��G��yym]W���`F4U�/)�"����E�6�3Af����s]CEt���o����a��Vv��c{���3׭ټ+���[m�ȏмu<a�:�hn��\�r+Z�V�.N0�gV]Q�l�SU�\�3���Ex^
Fq'$�O�"#���%�������(�ˮu(술u	�cƃ'Gs�!��omS�>��nxo:��\?PO�>�J�����?n��M���D	0ľ��?���^+�ኖn�� ��z�e� ����'b��Ҕpf�i�O���3Ѝth,�,�Z�n�*�\���i���vƵi�FJ�&x⛥�V�7�U�3�%w�	>�,�}[6"�a�ݺT����	dX�뫲lgi�0	OE��%��ڭ�
�h��R�Npp�(�yq�W�(�;�{�9H��w��o��z��#�����Jy}Op�e�Np/w�*�yˍ7�oֵ�����h��Ð�MՓJ^�2>H�q� ��QgYkn�N�`�R���.*P>Yt|����.�p/�:�@�ǩ�R7^t#�)����y7�s�$e�����ᬖ�s/���C	7����ϕ�Ϗ��?$?W\����i�f_�1H���EH���D�k�=$z�5T7";G��D	b<���Ii����-�ԐU��'^�Z����)%��7c�ؼ�mO }d�:����ONR��Q�Y}dݿ�5�I���\�4�,���GG ����w�,�Sו��s-�[�x�(��װz�)�a�3�'�]����X7}�t8�T��;=�e/�K�*�Vk�e���W���=�9g�֛:�ǻA	F���8S.�&����Db)-R���qem��B��l�@h��v�a|A(�A�.�u_�����W�ƨ��P%���^0�Xx�4��I�2Կ$��XBA�an��D�7�}�)Z�ř�^��!Y���� �a�n
ĀCzaߋj�1_os_��� B���lp9w�k��%i��~I8��p
Ư�l�=4������ƫWaؖ>+*N�h4�5쩉�G���DK�RwXO�&-B�dE�w��̯�EXÜ�b�D��x]v�x�:�I�^��c��D|�����Z���!��r '�B�&����"#R2��-��?1�D�x�@�f�"�ݳ4v��^��b+)W�@�l�e�i�ncN������GG[e���q��c\�|s�V`BPv4:j��	��]�H�՟�/lF*q�ZW��ww۴�'�C)ͯ^�'�~�����cL�Px��%�h��� p�A�S����k%vjS)�V�d��ު�h���LKyI\l�)��P̑��Q�f
�9$�*ܚA��9̀�}'�+غ7Ȳ�R�A�E�(z�7{��]�a:fwu9���~�o�{�Jz)	=Q�K��8�vC��Xۉ�CϤ+��Ѷ}ڵ�Mu%�n�:�=|�g��%k�9ٍՠ��+�$a(Y�5�I�E{�&�R�BB�\�W-� ��&���<s�?�n��Ό� (L'�XV��۰vژf�:;��1إ��a�X�=�ԯssb����HLf�u$d�۫�A�Z�|�T>E�_�CU6�+��,/�u��Q)�4X@���شt����0��4.�%�������|�)7R�ے��9tF�?�ʰ-)��-�-0��޸:}�l:tqŞ��K>"��=������ٕ%�ʆxy9����sO�Y��_S����͍p��|�I-�x^��hj��>�2ns\$_����VD\�fOJAӬ7�B����!\[Vz�������m��Y�|�%������ �/�s��I��}�m�$ֱ�<i��}
٤$E6J�Q�h�l��ʻ|jȝ����_�ΈD&z�`E×
��'.XT���n� O��zl%�O�g���kGז�:;T>�O[�n�^�%�D�W��r鉧\������l4�;A�
]Te���#^������%�p�鲈��i����)ܯ��}��Tٚx�3�PQ�����UQ5����Oo[��W���k�4��4(�QJۡ�:�\xc�3C�9�m�{UŖk�B0�,+�Ò}�s��W/�Ɣ�
F�ګ�m�;�(��R�"�U�S/Vp�.r���,}��B'J�vp�G�0�����F����O�&0&�e�����n�*����w���0�7WhKN++0Za��8�5��K+�hu<HE�k9x���-:���aK��I�7�h�4��7~hP�Y�<|�瓧�Į���h��)N]Ь��9�y �rl�x q�@����G�6S���c�� �P4p J�@ݕ�H��Zh�X�[��%8�E&����������R������ba8���a��0���,����0�w{�0���]���D��J���{�PD�(�;��M��aUN�/
)��*#�v__H�� �>��b��d?eB��LCy�Қ�Ro�Kq�����`=?�1�;�%����Gn��a!B�D�&�<�Y�!���A�$c����7�B��z���[���#�׃n��Lف�TO �(����`����>�D����Q��c�fꦖ�am!].z���/݁��p]�x!��aے��[���nB��wNij�z�ոQf4ukҽ��;�_@ �pt=(T�$�}1v�8��=�Ł���6����X<y�5�;��s��sk��\�4��R ����0��?�m�8����b����.�wh��־�ܦ:���Q�|���u�w�@�T���-�Y+K̛�|@(ƒ��_b�U��\��d�ȓ����L�og;+1,�̭U�n%#�u{���mƕQ�=A���s�C�� ܽ셌\��h�7h>�Un�/m���$%�r�
Q+�y/��������焃�NYp���G"C�p�%�.K�6`�}��γ��l�w�&��z_NЍ�V�&�,m|H�|�L�;V�]d]�x�-��1|BQ4�(%Wv�ixe�J��ͼO��A�
8"�v���;�PQbݜ;�'B�?4����c��'F��8�Z �p+ �)��؟�C��D�PsF������!�e�>7E�ٳ�EY�-�|��W��N��/�Y�������^��)�8 #��~~i7(<1B�JB4j�4YL��E�7�.Ie��A���~���qiƸ�M�i8�=~��:~��g���������x���������x&{c괘��X��mL�K!N�)��$eV�lVu�u�r��"����u���UQ���Z��0�,VN�P�� V,�!���#�*���E�����U��Ϲ�G�s�2n���c;� ��z�Q1Ʈ��A%Ef���O_��ܷDϝ�i$�Gv��f�f�t�;hނ^c���F��]���S�T�����3y�U��z�ʕ�e�k��05X��9�I�TrL�:yu�$I�L?�K�ep���'5��#�&��w����������=y�r:F�
-G��&������Ϭ�e���=
Ҳb�-��]Ob��W��Qf��m�� 5��;=�1+�ifQ��v�X�����(��-Q�mcJ�IqUx����.�$��m,ĊKg��:�勱�u4����S��C�WT6c����G�y��>�:�g���$�ƞ;�4���;�@Ó�k�`ߟ��q�8%DA:�E��V>��Y��Rhl���@I��?���wq�l�06z���3��ƙ��d{bf�x<��&%�>���R��fն�R_���Խ����g��'2�Ⴍ����� �������*���	_�S�B�﷠ �J�o�8p�!�Ԃ)T����N�˞�Huf��	5��L>q��`^�9�G��_ 
p����K���<��f�`��J9BPN�q�ͺ��)c�l��f����W����׆��[o4�Z�X8��aw>D��5y;��g ઙ�m�%J�h��9�m�����D��a���F�>&���$S�<hZ\�L�;^�<�W���@�U�� ୸͊`<�@��(���W���@:���C4+�XP�)�ޚ{E�PDW����s#�m��AW5c��t
�~1�ce�Ȗ�V	s-�������;��~���fE��$�Myf��SB�=�������v�씔4Ar��RJ�̚��!�X���7�pO{uU<�"�F�G�L8��^�m�<���$��
�����rP�+t�!�G?�R�B�W�DV����u@V׈𐕼x���1z|���^���x��O�˲ 9�]�dOz�|��������_�5�4l+�W2Y!�X~���J'QrA�2��?��U�J�cXhf\�����J�]3�f�M%���	�R1x�*��e���"����}�
����b��=�}�5�ۍ�RnA�tP�..�J'%�^ɪ�^�IX�˰��?s�Z_��ȓ����e�e(*�g�s%����B۔F���c����r�Q��R
���^���ʇ����.9$<q��%�#:ǺyW �-��Ds��$`��!}��h-$�컉ʗ,#�`��֮66�#���h����/�,s)��ħ��㝦���}r]4��cނS�#���������3�"��mi	�M�좇r����@r�/���ޕsј�	=��Z�h*-�XF��Z����-�y��G#��'-�n�-ʔ����%<��j��[�� �L$�� �#��z�C71��CK��BS��p�޾R��l(+E ����c���0��L�9	�(��0w�0	�ۯc��_�h���n�`6�[���`ٟO_>����<� ��O5~5n�}�3��;�9�U�q�+vLq��Kg�\���1{��w&W�$���ɭ�5��N���x{��/RI�_� ��
����?�z[�����W�~�b�T�NR�z�>��p0:�%y���h���Lh�"���@�¢�N���CЯ9E�^����/N�*�_�oq����@Q�oS�)�P�<<bۖ���yޱ#����넥OQH�]@w��o��+&�����s����.��N�5��W��;�%1�Ӿ���[�9Ye�'��'����b��PA\>�!�mbwC��x.M�L��8yvV�	�����*)P>�N�*�I�Ȍ���娸���I��oݛ�;E�)eE��}\�]����� �^ܢ��/�\��L7VD��j��t?p����;��_��XWMg�������!)��)���5�aĮ%�;u�F����,��s�r/�BC�ٴ;� �
*>�������H缍��Xx4]K
��2�H�"�#�UQ���S\%K��D�y��h�#����y+��E>�,��0w����R��>������"50����&F6�z���3_��zI��9˟ 4����r7��q�C����0���d�f����(������R��J?+G��m}$��J\]���8��C��h����(s��m�S!#�-�Ǯ��{�����2BA� �㟖��(��b�	����Q��H3+�����/�d�P�C��4��)���������2�3l�΀�,�������%5PH�j���7����}������[�m�ԲJ�|��5
�n��r �B���A2�Wj�*@��A1���և�9�i�Q:{~���P�꿚PyȺ�R�)��ԙV�ۈ
�_
�[������H����,v���{M�mI7R]���uYjK��~���F�%���4%(�6Z�C��@��ͫ�M?s�E[$v�ʂ�EM��*!��U}7�$\�J9��W�OkD9�_4��-k������Ë����&_����.�Կfz�I��D�].��y�.xa��[�p/�#�T����t�[m���Ѥ ��c�_��1�K1(����Ni�v�||�..��|�ZY"�K4�E�<�A!��Z����y4���ܬ�gyfe��{q�0L.Sq��)3�5,�?�S'D�;��g{�A�ͦ��B���\cJlz/�~��z�_��l���� Hce	��Q����? Nۗs)K_^Xk��.;���5���
�uVO�l� R������y8�9��)��T����5�t&�䐙?�D]%O9�5SZ�5.
�Sc5�����$d���	I�rTTmC���C���	���ިl�"-�	{��]���h����a(2��t�k7���j7U��X��;�8�w��ȽG������B�}�Y�@^V�B$�+ȗ�B��fPa�`.+gǞD��h&��p��M����;�@,��j4�ɏ-�2l6U@��4���A?q���xl�U�yK�X����y��m�͑&��p	#d��i�NJsm������;��*�/f��1�>+�7�q�=�lw}��Y�9����>F6jL�$U�'�
��t=�X��ן`$2���`������.�)�-��!���Jq�ܥ�P*tok�o��aB�
w��n�P�����m��م�}�E� �Q��ȎIE(�ŇV��f�9Z�|��!���]�e���b@������ Z��+L������ini�1�e$�����w@jԫv���y!Vo�߅4�-�l�$�b�B�����qa��r�=r������
Y��t���ɎҺ�@�ʞ8�\��r~�l	՗���} �䑶��+��l�\�bBF�w��lI|�OF�-��d{�u�W��v�kM+��*_�7�oS{ܵhR���K����y��Uv�O�
<����~����-���6	>��7ӧ���HW�d��댫q��V�=>��+E0�+M�aQH�t[��򐦘|,~m23*ڈG�x}���2��t]���ɢ2��F�:]S>G�q-��خ��%�?��B��ݮ٤�n���$�\V��a�%��ۊ�u�S"~�"|g�*Fmu=�b����%y�Y$=�\,_ :����ܑ�����(T8񂻆v�p�Ҏ�T���$L���/k��䔠��޹�	l�B<J��9�XS��rK|���H|[��������v�8�K�
}��������0(;A ��#�&
h/%���
K��Ŭ�$m�а�����2�����v(�}d �$6�����bz=l̎쀤��n_�B��/��H�k")���tN�� �
��^�a�' �5T����#T�+��*r,w���B��Q�?Pu�6��y�
fV��i�b\U��iOuGabY^0-�{��[�����Au���p{���g�#���uq���"�8$0�9C|��� ��K�<-�p�B�WU4�<�!aX�'�]|��s���P~�o�Qt������~+�����p.gZë����]V]�P+̆c��	�x��Arڮ���?���"��nM��K=^�1�)7hL4d���������W]T.A��A���!��4�����w����A�n�^7�����Z�亟�56��)����D)��E`̦-"�p��`WFc-��m�#�N��m�N���Lq��HUq��,�DeJl�y��ε����[9�3~#�K+a��<�1-���0#
d��oIY|�r�|��$Ȯʸ�I�*~�R'{2�CE���J��>.����f�W�7��i��C܃���~鰔3�{�پ�ǣ�Ē�����~#t�0�	� �.d�EAk^�=��Ǣ��x�q��g *I�d�8->@n���5���d�7�W�rm�s�?��鲌�Z3p�V�����-ePc�}�Ε�q�p}�5T�=�ݏ��g��z��;"�c�A��E0��$�Z��©�����-�D���g���;g��/�^T� ��}�! �����K-�;���Sħ�|gt�����LR��F�\0�P:�Мsq>;vg�� �AOC(�ZK��$��Z`1��d��ƫcc>�p	2��OI��%�Mnν3���Ӯ����	�I�vy��S�/�KY�l�q$�Cm�:����*��I���sӀ	_X�$)�ɇ�_Y�� `)p�e9j��4�>BU�)��O���,��3��.)�H�:�k��vӸ��T��S����řAdq���\��=�
^h&X:�hʕ���{5*-�o��<�*��L���/uX�
&0�C4������V��N@6��uǞ����Z����*B�.� >q�N
$�\�m�Di]���gN1N�r6%�nV�S�R���ϕR���ǧ��h`�`��h<����G_�	S������G�	4��m��9�C�HO��׃����L۠JV���2�R3.�Qf���CՓ�ԓ�Ud�W�'�$O�ͽ7֗��~��[�?B�N��VhΥ^'B&(RN,����F�U��LZ`�Ӎ$��Hә)��!��
��f�o���jn}c���o`��,^E�ʃ�0����W~�d�?
Z3���"����ʩ�(����^�̊=09�z��4��3��[^0��ͺڬ�`y�|�3��Y�)�2t����K{��i�pT��#������=�Ĩ�K����f��uB���T�D�c@�#05sH���ɧ�ގR~Pp�F�vね���,�q�sC�y��ifvD�^�C)��rc1�u��~rAQ�p ��2������7��K�w���Nie8M|*X�X�g�X[�m�
b,M�t�1Zw�K�}�9�	�G��;����tޫ���ՐsO�jy�M�-�T��`�f��"�I�5F��TH\��?������x��W���C!��f�b���^Ez��ʓ�c�Z��aZ����\<zC�vwrFJLwh�gC�{��G��h�.�5�stD��7�Ɍ�:�1�ܗ�`��)x��AH-�cQ�m"�
fBv�O���?f���n>C8@�*��=2p�H���Iw���B��e��?}B� �<𾺬����H�F���7#�tg~ٍYiHSd��7��ᓤ#�(<X��$4� bh=���{��a����O"���U��6�����>\���U�0��V�s��������>ʂ��U�����'>r�Z�B|q�Mϡ�>��h��Xk&Z<̡�37�G�ot' �A={�6�O�D��0TP�����%�_��+���������Z�0[���GȎQ`���'��D	@7��TT�ߦ;����*&`-u)'&�J.[qC2�@��sYyUU���L[�H�:�CM�,\�B$�Zo��ܝ�N��ߴ��0FV��	YB^u�HO��9W`x�:A�]GD	C������c�0%�#P��4__b�'�1N�����{ҝ�.��l��Oyn ��]��mԚx6�$�Jn�XJ�d�L�LoGW���tz'��n���c�����[�$MaH{k�s�kL�E������#��k��0~�\d����u�b&��uJtc��璺����Za��׊����œ*���� o�.�r�"��]�8�N�}��?�4.{�#�:�G��Y��V<%F�մ������r��6�I��j��-P���@�%.p�����Bm>��F�!)]}f~L��8�h�k�u��2�����!NĬSӯQ46�G�@��G�y�_���E�Ⳛ��g_��JLkU�-�eV�PSņFBm������M�&�i%:t*,'8�A��"�q�&�$䮬u"��J�WG�!s�L����kN���n��C�iR&��x��W�]�ZH�7�))������i�#N��{�h�H�C���M�'J�dZ^��&t0$4;�Uhm��+����(�]��BS�]z��㳌�Tݯ�/�6���jDp����'ę�5.Q|���1:cޥ����e#���xʅ��� ����� �\A";��^1�{�i���v��A㶰�;��2VuLr#o�k�����3x��Q�؛|v;|�E9���nZ4f��/m���I���!�хD�L��r��+�G��s��g4���w���a:�wk	�p�.��i�lL���yA���$	����t�o(A������p����1���W�vy�A.�mI-�(���Z=!eb�.�!��}VL�- ���g�P�K���)�֝^��*�󙴬E���W�iB���:�I�����w -e��|w)�D;S�ܺ���<V���I:88�j��n����u�[�3�=o.�-��f&�W�=qYZ(9�aϸ��z�ht�ϷDr�a�r��yB�#c�9��+@5�%���h���&�������pѾ-�.�%u�> 6�*G��IbY^U.:0�fW����OjX"=�'[��s�a�����r�p�TZd�tgA�P(Qҏs�i�y��A�������P���_�xXn��A*��r��Wd\i�\v�Y��3c��T�m���0�����zJ�D�󠠹���#�����ɗWok�Ebi��p��v�j[#�j�[���y�����XZ���r���v��I�{�S!�����]�/}ϒ7��P�҆�ֶe>{��_�mɐ���ٴ�aJ.$�rF�I�_�Ro���(��X�k�dvuT�4X��vӻ,[���؂��� �=����Rȉ��/�	�J���?�b�\�n~ �@�b6�B2�1�'�s�tZ*t�4����#H<kKZ�,��[�{p���m{m�>9�u5\�5N�&O���C[fQͬ�vW''�9���W���S���h�+|�b3�Z��Ag�d])v&���Ql��Y�j·�]Af�A%9MT#�ס����L��هK�N���-ٿ��1N�?e�;���پ�µ�i��ZJ((�/(%�?��f�X����-�.Xk
�'�U�l~�ȸnj�W�B�wB]8�����ukn9�&�{���h77!�`�vW�ns�K�s�[ub@�����wR�\+��T��'-{1J��/)@ϒ�V���m���nq�r��.��!�����i�d�m���������:Q��MD�w���=R�<�{�mq<~0jb4����'Z��@�G��P�-�C��jV
ZB���:mR�x�m5h�Ѭ���������Һ\Z��U���I��!�&jk�D�$Οk�˻9a�'!B����U�P�E���9��;��˄;@��V&R�O=��Ў"Lp�����"��oX�������yɰ��4w�R�`P?=) �<��N�ixZ�V�]z���:��b��@��N�zAԍb.8��P�/�>ٕ�3R�Ԅ���GaV�Ѭ�A�%U����*|'���X��NY,s{��EL�_c��+D�2���˞��s"�� ����8e�q��G+����sL^�]��DA���p߁J��x��xy���1� y�E��P�nY= ٔ�T�	hlj���d��c��G��Į�.���q��6@%�X�ȇ?��9��q"�es�����@x�Ai@�"���F
�w�=�$��4�=���'=;��~H3py�U�p=���:2˩w�7Ļ�T�h�����}4ђ��v���Z� �yb���di�ƽ���#ɖ���2D��FX�	i��dP��߫���1�bR�����_rӀ�� �S�ai�����q�I���Mq�������^澑&m|�DFE���6�N�'uFB~zf��F�]~K�~�d"�+y���D���Ę�%��r� Q�w ��&ޣj�a���}�O�=t�\w&�������WIB��N*9���ʥq޿w�1�@�!��5��z���Fk�dC�����{*zE ���ӹ{ۦ�ƃ��Ie��� T��Ie��Y��\|��>.�^K�ԎW"y�����g����	���/ḑ�^�W�9�el���q�pS�<��_ٶ���fFDQ���ў�W��rؔl6�ឲ%��{���i�|�:���%�Y��ppCp/��7E��*pI*q5�	E6�� !�}����bt�9�i���>�7s����1�����! ��Y�?N�b�"Inq-�v]���}�p$1?���/N{�39�k&-Í��t��4�Jy��]d�/��/��2����G^��9�J������];���0��Z���f���՞��{�$�Ic��p��,<}���?�DR aZX;���� 
���SX���k#�c�F�aʡ�JiT~���� $0���B`̕�-����s�:T�U�8�XVWU@D����5&�T���d}^�wm��/g�5"�:!:`��u��9Zc!�u%����_�P��DJ#c\W�H�#�I!'����`���B���);���)���J��[u�e˶�,F��ǭijqdX��\l�]�;v5��^@ɏJ��3d�*��,tCDg�8r����a[��n2��2�C��y3�����@f5�|CW��t}D�����-nȍd׽�i�E=���"�~����P�ڬy��A~NH���/Λ����W�b�j�T��c��7{_?��"�l