��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1eO.�l6�?,���C��Y�S���/Fka:qsF�4����ϳ
�'?h�^l��yi��g�^���9��(£�dHB�Ȉ^2���\�"me�w_���80�Վ}��y���N�[L3q�\\�_�������D�<vhy��<d��ȰuM��Eɏi�c�3�꒑V��XQ��땩WW��ݽ$�)5(�s��ZO��Q���8��7�5��u��V�|P���98���lGX����D�xIK��J��s`�x`���4E��@��>x���v���.���%�Z'���k3�عӻ����W)���� ��UA��|^�F�Ҭx�}���V��E�-��q�yP^�E�1�:a�jae,~�]���A�P��Q��A���NPl�ދ8�bIə��G�'�2v6�/n���P6���<�}h��H�P�%�E?"���(�T=h��^��{}Y�+���|T��zk���!��W��Z����@���9dF}L*9Z�:�ڿ�'��qjC�;����I"�����#@��r���)EE����a36<�B�J"W5�W��6	�y0Y1�a�����t�i2�J��u���T�RY&1ݵJiǭD6z�a����9��8��2N�_纊��ڂ������VV���g�v�sİ�0�z�*�/�>Ē��c�g7�}wm�
�
D� L��눖�������i@�}�� �6������ ��q<R�ؗL	a���?��A�>(~v1 x*Q�K����G��HsQ�l[ɻ{�U����"%?m!�`�m��hY+��1��,�[Pt�$[��Jȶ�x�Izbs%n������>�Df�@]kou��Ia�vL��xU&�C)�ΤniZA�,��*s�&r0ϕɟћN4��|��X}���sz�g��~M�PK5?�Z��<����M�h��^�d9W ����=7��g[�|�?N�z�)�;6��u�ݩ �r���>��-���|�´$�hr��`�� �����p��]s
�;(�ީ[�
kEy�:�\h纆���tb�K ^��ั(sg`�&�;�k�1o@�k!>qޏok�9ʰ�F����|\F�#�Ge��s�I�>mf�-�
���7��R��ֿ
�����^ =L���?���wB���Q�,���r��\S�5*�0��C.R>�Hrt��E��GI�v/��j���:�A��I��=�m)4��d�o�ˡ��k��d�Ӟ�\?�D>N��_1��1$o��vyl�^��q-h���P�Z򌻊��!�������l�U�9X��H�2�^�8W��+4�
\i!�\
�����սg��Qќ1��拏�A"uK/�Y!=�P��?j����R��A�ט�e�ɽ�Ѣ�P��y:�la(�$�8��y���s�j�b�<�8�Rr(�B��-���Sx��N�����\/= �is��H���f@�e�#Rש��I��,�ce�Nl�;��[��5�02[�EKw�Σ'薂`DcV��nք2�e��u�.�&��i���gB�8}��?5>�=�B���KV9�Ŷr
�snu�bxR�g�b�ԯ��Z�1����v����
D���@��ێG�B�M�������^q��Ȗ�]��?tv����P�|x�Bh�g�JC��v�l�f���E"1��+,GΎ)�Uq��`kf�5�b��Ff�ס����p^���W��<آ�7
e�c!� yK�K�6`�i������k"��qJ>��N������3|����h��^����g�17����},ヰ|9�s�o��2z����l��i�4�.!�<ݼ6���k�+�p���^�n�{����5�qNl��Z�sX@k%7pedҤ�lm"���)��ҫw�ó -}��;���c��T;��Ը0��8�໕Q�l|Mv�]6$�X��o�{��J&#�O���[���"'��̷`[���L�K�V��6S[��e�\?J�p�>����M�ȠbF��eX�R>���1����9-`C�
�W���j����!GS�`��"��Hұ�^Z�e_��Q#$6��ͷ�����E��¸�B,;��������)�7u���b�� *�	CV�>��E�=m�w>��A!��d��_���Ϭ+��M�׿DE �����M%%B�ֵq�ZQi�no����]'�2���Y4�<�%�W9(2�&=g��|�<�o�j�ۑNi���\T�����<�X>�ƞ�2�]1���X�6�k����H�1��@��5)�޺#
#f	�OD�_�T��?[~�]��d+���A(ޗw��dig\���2�Z�])��e�}㾞���3�v�%���=��� 9C�j�9'M�(�^����wG�j��^[�<�]�O��Y�����n!�;���ʣ�.�S�+5���D2U�&łܣcx���%��\���(m�a+���,�:����Uj5ґ��~��ؒ�����W_C���S�i��?�	�reդ������]��{^�0�O���;���������y	��\�Bt��ǣ�~�o��Q��&��X��`�4oo��oՙ�V��#�]3\NhV�ge��⯇��_f�KS�^��~>lfs��,\z�%�7r�U�zO�5Ā�{���40\�PZhG�I��4YB!Xd'4~��յ���E|ҳ�鵉��� �~1R�U����ыۆ��+<�{*��N�K���|&g ��J?a��L��O����\.�����?1rܔ@�,j,u
<�⫷�w'����	XĂ>��M	)�q�É`�:oY��m��*��3l�2�b�,d��^/�z�`��^��o�au��"�yl4Ս��(s��v@˕ն��kS��j������X��U��1e�~��쭑���I��	߫�}i�9�;F�!@ڄ�j�~��!I!졺�����$�ܼ	4A�j^]kαԪ������m7�m����٣�y$&:�٩�4�;CDCash~1�Jm���mk�܍z*�n�L�,����@>������T�ѭ�W3�h[�ec��
������t�jxK^ݘ�������q浶��.��[�Oik�����̿l�%��#�[F�8�v�τ��6,j�Zr�O�Ю݁�/gcK�t��#���^#K�Y�]�Ё�� o xX�۷,��-��I<=�g�nzv�Yx�(�mh�Jæ�+Q�r11g� �������r�s�tp�Dj���q�C�� �d�5���P�lɇ�J����gp���s3��G�X.��!$Q*N�j6�>:i�������)�`�@9�b�A��t�T֊��V+��t�w��~�.=�s�j�^�UQ���Q�x�hZ\����N��y��
�������MJ'�3�On��h~m����� �0UD��ӳ��jU��]8H"���M\Bt��CU��I԰��q��^ϒ�O���.��\q�q0�z����Oޘ�|�R�h�ϥRf��6C<��<j�8��ըS%S����!}��i�3�� �<fa���`�_C�t��`�;���w��bQ�=��"�Ig��Y�m6��ڡ����-	�� ?_��_�1KH-/�\��5�D�R� ��J)k�S{�A
�j:���w>���<T�O�6�tY���p���Z���.���9;�ͮ��;�F�K�&�+}�%~ =���7����:eL�P
��+ M�g��{㗨���L�R�%S��I	tQe��t�fF�E!a�__�P��t�ߓ�[d=+�70{�3j.��N~��5��qhܝ(h��;[�H��j�����8G����n� ��V��;�1F����l��LK���(P�y	���Ov��׌�t/Sr���5���rE$<�<|F���'!1.�ԅ�?C����E��b{lr`gƖ|�5��-�>�b���pj,;E�O�
bUͥM-���<�a���Ve���j`�n�����?�v�(���-v��F�E��iy��E���i
��Y�=��T�e�FN���NOw"{�g�v�:��кz���!���f����&��Ծ�$7Ie��G�(�q� �/��Ƥ�Flh�0��cIτ�kz���W�|�FLcg*_g�-`����j�Ͻ�  �-���j�ڰך�FD�5�Y�6��	�=9=������b1N��,���K5��w#Iiխ��V�N�؟�����+L;^eg��1��X���r5��bc�+S��M�k�ٸg|s����]�}�k8��l���0}' �=��(���<��M�d����!�MnJ�Q�_����v�Ԡ���Z!B�c��A��6��@�*~�m����(��y���07��5�k����HE�'����C!Y�S�\j���ڗJ�_��*/%l%�^W����*C,Ur˳v7�u���.vՃ�Z���K(�,��!]㠚읉bA�UB�ǗbD���of[��[�3ak���k��Ee��`66V�j�h����_�M�EJ&{��bs�a�n_��:"��j�B=���k\M1Q�3���������hҬ��moB���t�pV8��f�=�AJS�����er�e#�i����+	����{�*+��� g�Z�8ԭ�jbW�^x>W��M���u8}(X��Rק�H�� ,��J	�'�'���\گ�ț#��WcI�k��l���|ٴD��H������l,�zuc��9YWf��e8����B+��=��a�:Q��nZ��9vz�����]��0���t�����Fu�6mag}�H���[��4��+�|�pPop1](���O��?y2	EM`��a�΁2�D�����M;���a�r	�?��,Kmj�$
�.��1�p���!p[�ԅ&�������5Ⱥ��c	ɵB�;���<�P,mb���7��Ws5Sg4�9�|�qڗ�]"z�8v�w�s�K��i(U'q���ڤ�����;�+ȣmJV6��X�tr�ɐ��mm���c6l�!�K�]4wO?����坯�%�㗑�<�
�rE��>�J�mŤ�-��*@u5�"�[���0�g0+�ڌt1�ك�LTp���ּ�肂�͕���A��T,=�e^�r����x�L���ȵV� B�pE���׾��l�:
�����5�e�7�)���c�o���]����k�D˪�;� ����W�!XD˗�X0����h�>��y�c�o��Z#8-����_���Z�~x�~�Z���YN���ʳ3Ao2��'%=
sDtr�dc@	Pz�}�P�l��J�s�?{<�-S[h��WA��k��[�"�Ϗ>l�+�>��¾*�Ytx,ǁ!�AvU�w�"E�	<��)�K�@������>��Cc�M�6�]�{���z%�^#�T-�����r`l��r�����eg�J�!�L��:G���Nr�"g�?�:��Ƙ5�4������"��OY�J&��.v4���4���y�Wi���F��>Nl6��/J�X�B#��uh��Ƥ�wI;�SB��l�f�_�kg�X�~:���� ��V�E�j?�'}+���#���m)���l�Ϣw�m�7D�6��L�Ւ�z������C�)��造L+$�Q�(3�m3Y:�G��-��Q}��!��k��TK�ruX~��;4`';X�Ɉ�n	�Wj&g֜���r�l�V�pdz�.w�|��ܭ�N~v����gI�l
��.3���r��1����jX����k��.��Q��S�	Yj��ei3��c����M��$C���u*ܬ�2S���D$��]�}F�N�+�Yvh����֓�ǫ�-O\ H�#�x�������$È���X�(�\%X��"A��Qb\~9�QӋL�4��g���1|֋9#0(�b5g��h�M��%j.#4��7��,PL�o�V�E�*P}"�1M�����`+2��U���ꔓ]g^�?��KC��ʧ��?C��i��5�:;y������9����-2sy`���_ s��]���&�~3S��M�Y c`���0��W|{��;���/d�*Á��d�A��ñ�Z�'�K9Ȗ+�0L���&T\N�t�����M�:Ѭ�w/�Wg�`��74��d�H�0������8c�6�.;�0�����X��*ɳ�7������3J<�����٘�·���/�PEI+%=ф���3`��j=�ԑ�)��耽�:m!Mvs;���k��pҟ�ыB��,H�d�H��)�鐩�f��qN��8/G|�"02�Z�o���=��u�\���]�2�O���9i���Re2B�"���ed���}��9���TF�(C���|��E�r���Q
�*���!�i��;!��	�n�u<�"�z�o��� ���2I��@��N
|�q��#���h�Ⱦ.v$
Sv�YI�6*��ʦ���]�]JO�.C>w��_%!�a�1^/{�W ���f���Dk�Bm�~���=BV`W( �5��,�t��&@���g�
�i�T������45()&��ɨ��U�S�b���~tu
sW9��fI%L���ǋ���Y���8c
W�We������E�� �Iꀶ���]�.l�����[;��On�L��Y�4���(�+��b� ���n�Z�ۉ����B����t���,�W~�(8�A�Q<"�Ru��-|QSMc�����3���t|��'*��n�h3U�l4��!�,��CF vcO�w�R���4+a!�`�͚5�@PB��a{�ي��t��0���v��ޥ���ȌzW>�g���2�e����3˛��x�$(���`�A�A͹�b4AHA�Z��N޹N���wm}��U�Y��2n#M�X�!�����a�D I��O>k�d"+ȟ�cU
�'��A<ԏ�e�@���4P^E#]�-;8ֺ�Y�q��:�[3�"���p����g��{H�)O}H� K��۷`�{5����G��(BN{���s��H$����o����!���� �޹������n�T��n�5xb�gd�F��m�&�eS���r�=X�:��p	w1�6�%.�(=��Z����w>+Ղ<��[�o�Ť��(U�eG�xWć��pWOX_,z���EI(��b�S5�D�)r-�rUTQ�M��?�.��@V��'ul�5�Xl`�p1�Ň��0Fi\�Ak�&���GW�2pOu��ѿ{L��@��Q.�w���ͬX�5�/3��:�t��ޘ�{x��7C3c&�~�4)u�S�p����ի�Fzs��P�Y�*�~�0���λH6G��'N�^�K���wg�&P��|���:U��ݕKpR�8ϒv�v�����;��K;�|�H���Җ�/#�����,P"Ѣ��O�Ȉ�e��r��f�W����<g!�63��V֞��z��������y���-���MCG7�=�v�`���ґ��]����:�e��p�;�U.Р�3�1ů�kj��MU�O̓�АU4�*S�X�\Q*�����g2����´��;쓹zTFK�����0���I��ً���Din�C�WFO&!)�� ��A���I���<`%Y����h�N<��W���bpƋ��x7֯�Oi�٬#�}�$~YL-�wD�;���GW'$����>^Z����3�P�d�b����Cdk�v�a��#��H�9רq�Lю�G�q� + �r�G?��<�|�x�C!	�Ӝ1��/v�X?��g)5��k��%U��2e�oMB���W���HMW6����������Jyit���C��\?���(h�:i{�\��\��Ԏp��p����Oi�$g��4]���!忐�s��{�7f��Y}��i��GqĦ�b�w	;��u,~H�pn�#�����$3y:#k�� ���:}bL�;��H�(��G���P���*ס����{�&�LW�N�����q����.��� k�A�B���Il�.�j��Xu���;,v��E!�".6���:�FOpo�����#v���55��'+�G�F{Ee�BF�|��.�7;�#�].q�8-���hg��7U�&������? #<U�e�zzM�U��(��PGU &^h]>"3Y�U�P��o�nf�g8S���w��,��z��Vr�X��`�����/���w��?�spC��"�֭%�\7����R��*C�y��B��+�%��5��T8ﯔ>������/�y0���h��$n�A�*'�>�3e���/SE����7���x����GuԤW�������{�zuŭC����d\�I��,
K�Y;�?���nF�x*k�{H^��a���S3��!�j8�� �����i��?8�������?[�pI��M�?|v:͋��6�d�2�"G�6�c�^��*H�w��؛H7�	��cD�q�����M����OJ\C$���)�3�o��a\d�]Qē���]v�ۦ�<@�g }v/�q�9��V���N�ؓ�pOL7��U�M��p�����9�R���R����,�@��ܞӨ?`�/ń�1�VI��BFzMw,��$�$��l��d)&<X<x6p�&�v�c0_:�r'���O(�Ր:n�7���ęl
9	iD`���
��;�l���T
�8�Qǹ��!/����hǂ����ͨ���}��C���qH�<�	�:jA�Mhױ/+��d&i0Q��?fsi�Ya�c�LۏH2��h߆�\�-O��ܩ�!T�e�!���ȸ&��`�J�gLy���2�>ˆ�$t����k3����+P]n�D��sM���\������()}!�h��ٱBA���82�:���(�k#�=�)���zg�),Cu�w*�y�lsR���N�#����8��!��boDj�����hb��*�3?�"Q�?�ax��8#��`":o��q��xݟ=1�bT�D�JY��*�қ��I0Y�?ν�@O�x�Z7��㳔	��ݨ�tzZ�\�ܜ}˻Ʌ9Y �X���|��9@a�ḏS�k�_J�� ��籠Qhx閊\% 
������>�b��G�9�I훐+��v��� ��"�t��x���o�s���1�k/��:D`I��0��A\��lP�<l��3�̋,���
4�(oM�O�c�?>o!#.�A�4/b�S�3B��*�w.�BU	V$�Tf�/��9�,��?��*���e)}�{K�xOnBr͌�����Ն��":R�*��/Xdq8˕��6�B8�����)�q����O��C��h	u��M�gk��������UwY/�`��!h��\ο�k9�m➷.nz,�^)�L��~m�[C�|_����<�0����Z��5�4av5|���E�^����Q��U����Ƭ1a�+����/c^��
���������UN�D�Z��'Fm���zy����]JP�1	 X�<�(�{.7��i�]��Iv��"Ƿ��a� ����͇���$��J� G���X�v�Is�����MH��wڜ7-ڛ��[gx��h�0#�|^YS���Wt�p��L�W������cC��8��}Fj��d�2�D��d�D��!���+�r��G�W��F�k4�锵P�����	���T ��Tzu�u�hrcQ����AZ*�`��ܨ�4�6Y������Q��a6��<C��t#3H���W�p�]0�c�n��vp`��[���%:?�PϐsĔ���b,��E<���Öb�p����{,]O@����BS	Zg��&���B ��?e.��7'<Ю`�O8Ȟ���vlge�\gb���6�bu�-!�CIB�Z�f��^Q�Ty�VY>x�r-���J�B b� ��N��@��nU �<�����^�p��
�g���F�u���=��I6�^���>I��^KV���d�EܱJaBs�\�D:G�+?�|�A_�jza}7q˘-�HiPw��%A���>Sl5k�ޝ�Κ���D�ϊ� �s�7{ܗ���2�e֪����MϿ�Z=gq˩�Q� ��!����<LA-4���X���Y���-l%��Ќµ,�1�����b�KxjGP�iG?�Ǘxh�'s��\��L�0!���2�wHCD���x�TZ�^?FӅ�LvO���!ۇ���j�i��Jr��%��� ���w�y��/�OE�ߦ���}���
�l6�dJ+ֺp��0���U"aACo͙e�,!bM�5��tT�C�d�8ʹ&�9�i��+�V]{����h`����(;��<�y��yF��Em�3P��H&.�6��i��Ӎ�`pt�l#d	�!��W�"�AH~$X��#�^u������$��3Vkb[�� 4h��:*�&^E`���QL#	ůz�C�Y&��L�}���a٩�J2�����|F<��L$��_��FV_	:��r��'�8�y�!�0?�`� ]�ρ΃c5ֆ�J%.�L�Bz<Q��L<y�)�{}������Fzw �HT���2�9q��:"Ci�2_�&��B�xK6�AZ�,C���E����?H��"1�$�_���ģ՛��U����O2Pg���0/���1/�Ge�'kcҜ�A���?�F:�={����r�"mnl
Uj���/���0,rpDf���EɁy|I���5���	y�"j��3GQ��8�ߛѴ�fWd������R������F�'�i���t$֋tă�/>����+�g���H5g����U8��)Tw<��B��"ÀB/���ij<�a�1U@%h̎�抶9���$���#���t���cn�ߵ� ,G�)�|d[��G��?�Ͻ���׎�i�rLu�xxgظe���