��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��E#�1O�^/Ĉt0���0'�H��~;�.'}�;"av�Ux���r,�*�������_]ZQ��f�9V�kU�!y͚I������8q�G0,���z�������n�4�c��5��62�䗏���;�D��9V���}�$��|&؅�&�D�8e�����`�����������M�V���[��u����?���Z����o0�We����;&፟	�Aw]>�g-��_t|�k�T��sU���S�c㟣6�9I��v1^��N��(Tf�����߸�	�D�l	D���d\s�oX���Kq�3�Bq�qW�q^	/�]=�h!�i���\d��*�[B0r��0d�8����$�)	�(��a�qGwS0]x�K�Mo�U<2q������>40�̸
o���,��A��#�d�6hu���̰�@��+��EL'k� :��.�X���S�IgK��fH"]�*r���u����?����c����x�>
��	��݂�YM�^yp��j���"���r��Wm0*�o��B���?�<5�b�Z>�0:�C=�V�,Ր�-�v��VfPF�N�(TN��>��Y�|+�	}���`�$��@�	����bP����8��S������;#řE��I��b�̬00����BG�9zSb����H���[�+9�ϊ0vY��"�4%*S��@Y[�S����>�|���q�fk��*�����|�ՠw��`!�T�F�|��n�wN�o������Z{��uP�Vo��-݉����I����^U����fq�&�Cscr��!UY����2��5C�k��_<��+��VÕu�����GZ;#б��TM�"`��y��h�k���Et����S�}u�r3�rS��sa;²,�XF���e�H�d`^�%�Hs��w��x;���q$�b����=S����:<r��qP�C�n̻%<6�ڬ�����O;�ۣI�؄�>$]�@���m�t;�㍈}֧\����[�0!)*t���X�K:,	��H/~�Z�����E�T;�q��LM� -4����;�0�Ӊ"��|���L䮛[�p�ژ��� � >�e8���`o�f+'q� �)|Ĝ+��O����-��^�O�y�ݣ�B<j/�7�iJ���'�Y8I�P@V�ؚ��8�nU�.%��@�'�����E���66�v���w���s����ݞ�Xk��t�!�O���{ﲆ�[�|�ӳ��!f�"�� y�x��1��QS�$`��o��%p���Z�^� L8m�$�8�^1�h'�=���7�L��C?�[x�����w�q�o%��>�I���"�:�N�=����図� ���+�0�2u?��*�ܥR7�^W%H��}��s&����qb�ר��@)�k{ Mŋ� )P����]ZF]���ڀ����H����FL�咿�U�=:�W�p��̟=�m��m����~���iEX)i��kD+�5�Յ�9� �<8�F�����M)����IG��z��'�T��W�x�A�`p����u�@�\V����O�jT�-�W���&���ǩ��z�Wzg�����a��Qbl��`I� �:���
1K=ʒoJ�]��+r|����z��%|&D�4Q����ƿYd-P�Kw1(����073o(�W��tX�{��՛T�o��*���R��N%��t��^y�R�N�T�ߺ�b>��$�荐!nCX�c�N��zIt\�����o�)��|b�j���9�z�J(�:��ɯC��g�9ɏ��kE�y�Aw�3��1���zŠ���倶�҆�X6&K�Ի�"��.�U����۶4���	��J�n�3�Ɵ�K�6��	n��ۼ�y�i�3#�����i�a釠��Rq�HL+�;������ǁ�+�T��� �{Iی:���ii��Z!>�?F��=
�~Š�
���Y�55�pR@Q�a�i��,)[V}��l�lZ_����*��j��S��î'V��G�qA��td�`g��6oҽ��k�.ņ�@[�SIix��4��������ƴר쬔�����~a��BQ%6LS��K����~+E�qI.����_'�!��d�f�0�ܘ!90�U��w�	��r.�Y3���Υ9Q�U=������T������YH���gEz�À�a!�J0��&9�%"��y�>[�Ѯ,��Ï��g3s	���tvR��V��p��qޔ	��K����q�{W�!i�F�p�<�R4����QxhF_,5 ��ߐh�c0���>��p�ڧ�2�)�W�-]욞X�3�>�
[��4 �3�'VP�p�����z~y[_��ODPg,ʬ��i�zli��쩝�(s��.D��Q|��wQ�ί$��s����UB�5QP7�@�3�+�7�`ls'���b�����na�.�=J�gK�N)1?�80q�\b�H�z���u���4�au;�v��}�$
���t�|Ol��>7�g����^C��7�ܚ��@E�*un�X:���9��9�U�FIOd�I���6qq2,�[�m"��xԑ�pP�z���J�W�Bl�]ڍ*�"���5'c����Z�Z�&���k�yUP�b�e\wD�ʓ�U�����;�f�\�H&�{R R�/.�g��/�h�6�)	$.'q�Ҿ����!�Ɩ�a���GzY�v̻��}-U9�c�w}0}�����B�����IV�	����s}��}����ՆO�q}��@~>���y�o��(���m� (ʱ��G�Wx����M6/�Vc�L,a8��W_��9���3�`�^P&0@["��6]<���D.oB�?Ut<�0��U���o�W�t�U�fNj̐���M�xG�m~�Q����fq ���N��]�#�<�"lg�X@_R،�SD!�n3R�Ui�!M r�{<��eL��Y#H2.o?Mp�MR��ݢTQ���>�x�'\hK�
�"����	k��SZ.|U:�p�����+m������W��[g�0�c�%[oeA=Y�`~�N,^ P�{E�����p�{5���:�����N�K�վ�%uA�9��{1�� ������M_Y��,?��!�O|�92�4/���Y-BVS�O�üte����7�o�N �[�@N{�S].ȍ*{V��z���z�dYp��'j�ͤ�L�l٢�B�Y�Y�!JSg8�|7�8 �O9����e˘>2<\}�{DV1jЍ�a���l87�F}uԟ��Dt4�b���uuCo~���$�pg�3��T |�o���k���H�E�պ��xq��|d�Q	fMX����ՆAa��b�#� �w�8�7�Nq��U��<��)T��y�"�"�\0�_�YP��AiꘕC���b��!�v:S~}�� ���/�8���m,-�%Vk��\�TU��H��	���Cf֙��PJ�nՕHN��t-m�!�e�M�֞���Iܠ����ܳ���m�����4b�QE��&��n^�o��4�á���U��/b�OMA߽:jyC!̆ˢx����C&�0�x���![�BUs�ǉQ���R��o����>[O�5���9���FG�h���Oa�+G,6 �����	�܌�+���Q+�p���E�}Pq�HߍĤ.���/�%��_{�|E�MN�Wq�"��� lb�Uύ��X�'=~�ԣ5�hfK�揧v�^]˰�����*�q$e��Q����1��_7��$x�;����v�;4'�	��Fa�n#��O�� 1B����$���7Gt~�<��C��P�����J�7B�t,�-�!��M�@���~�Fɨ��	��N���-�U�+�Q '���������e��|	��k-����)]��nD�:�+j�Q�.��?ܨ�+K_\H�d��r�I���� �-�?�'��A6�g^4K;_7��[J�?���Wtp�R�t�%=���I��=9�R ��4��i;�X);d���_�8Cuo�Y���j�Z�}��"�MBM�j�B�
��3F	�S��Z���|��D1?�h�|3y1G�j��%�O�i��_O��6
��?�u�G^}�d��1�q���g�p��<�v�*�֩k��z�x������G-���]qo͛7vq��Ȱ�|I�N��e�J7#}�YՌ	��`)�{ĝ�? (�9C��� ��.*!�м�;�~�ɪ��>2��R�Sd�/;��`Z{�d?Yr�þRG:ڗ�~ro�d]�V.�E�������ϸ
ڳu�F+�KLVثDR�:�H��l�I>�G�ȕ}�b�����L��;,�.}�,O�R�ަK71�C�JB���.��$�|0�)�By�}F��
��B�3���$-��~�K�ȓb���rt��^�P`���F��C'�D���{�ȧt��䮕���1��:��~?u��NE�b�.��^�7�P�qp��dt�7��L�5���	ڽS���?���h���\�dZ轷�.�]b��h��0j��(9�Fw<��\�k-���O��fR�oA<T��;�4������é�����_����eteDR6�YWu\F����Q� ԤXZ�7�gS���n��mJ��6MBe(��E���8�2PN#)�'��Q�����!��MkD;b�!G��n!�>�J
 �Q,I+�)�Y�kQ��]	y��j�W�-l�`�F�T�8��q����:��PcH��f��@*o��wp��H\HR�'�/7nĳ}��.�9��� 4M�����4��RHm8���=ט���@�� ��u��܁TG��ϧs��	�ukF��H	�ur��`��$��W�����?�;l�{�>��<GB�!���p�<\��R�9 �*��s���cn��{	Z���@���?�w��<t�m��r�a[T��D�1�^;8�Ծ�#��)x��/Y�@���6D�PDQǑ�53�?2�\�1&>�A�\�n��IM �/f�9�H�>�
�e� ���]~�E/0�SI���F�fG�H�
�@Ҡ�	O�ɨi�|PfWS���[�o K��n�ډ6�+P`r%/�N��\W8�I�s��O��օD޲����Բ`>�#鶵���vB�ZK�wÒ�Ki�n�=������4�^C��j&���U�U�,�Zy�'WsP@��؂o����K��}�I|>�Y��ND�H%⢍r�/9����hI���V9�T�%��ao��#e��#�^"������mRo>Z1l�T}.=9�<���C���X�[���;��E7�^)ܘ���;�|�
oc��RY�n�I0��z��*�*�~��5\Yw��.T e�Ö��9�:iT�X�D�-�Դu(Z0�.��!m��zp�W�?:��hk0��ft ľ�3:u� ��^�#�H���X�I0@yù�<�mf$z2�舰�n��E�^���@�ܲ�zq�#��7W�3�s�V;*�J�T�����B��i�H�Ǟnꮺ��0yIz�"!z��A����A�J�`�<�u�1m��~"ʄ)32��4�'���J��k@>>��>]�Xbiw7Dp�ʢ��`���Y��]��uC��ja�2�M�?�H����'_$�._sf� ?r翛�
��G+<��Eݯ&n�ʾ�'���a�x��kQ ����GÄ�M���LdIދd�<��H���~)Y�	9��ҽ��U�>@�sZ������|��"�{!^��B��e�@��� ����g዆j�Z,��vʱz�7�9�<���2��\j�m���>�䌏��h�:�tQ���nu�/����d}�+	��Ԭ�q��7��qc��͈1�^R��qK��!6��p6f�Z��<��Z�7LƐ)�|s�#�UU8�k6���p�����$;v��� Q8�l�j�5�K�;�J�HW����3��lJ�:�%
w�}`�>��愤�iQb$Lz�����]%3�4La��I���G|�F�[cG�\=\ ܬ�L��g�����+s�dxI�!
�JP��My��KMϗ������E�}�sb^7O�tp	
����n9�؅�.�&1����V�ç?\�|IX��k��X%��h�̤L5��L���Ͻ�8ں#L"�^(���� �o��>�h�T��Z\�-���KZ{֧�RоǾ����i�ѳ,��
.��Ȱ��P��M�Y�}QY��!�_.�i�a�:[	G�57�Fx:� �~Q��o_w��Tg%��Y��M�.\��ra�௕Lz��/���4�1���#���\�d�m����1�J�T���^�+=2��U��N�����9�^�G��x.��CY�,��YT"
zvr�R�����u�X�~~��v�&3D�K6�<���7	�,��4�4oR_Z��aQ��m`����V,��
x�Bp�����8�l�mzN�s�s�jZ���쵪݅-�)%�/����f*��P��3Y��a�ə"�A���5�,3��a��մ��[��6_��%�âp��h�M3�n��)�$��֌GsG�bh�/��ymd{	���ഓ���yp�yO����[UZ���PF��O�d:�)#�wiO�B,���� f��=�xSd/S�_���\�u�k^c�=;����L1����c��H��e�Lf��cH*��n`�nk,�@Z�a��-�Ѽ��\ȯ��hE���ݨ,S���\����2ָ�cu�k8=��ޕSi}�NM1��kt�=)g/��U�-��N:K�>���
�<{���*�Zʾ��� ��Z�X��/�,�o$W{IJ�կ�{t ��j���φ�,9
uk�G�_E�6H��)�(.�m
�����^$��w���W�Pg[qb1�c��sx;|Y�R˓���N��e�mF��M��F����ԹA@<^��_E�<5�߲���?-�Qb��m�. �K��a�9AG�%�-�eƮ1t�6Wo	�x�i�{�i�&dKX��GǩMO�<$�g(Y�8�:�A&Z� A2�|Ř�B=���H�:�I����q���6��VAu�v�7V��}O�8��l-c`aJ5�����ËA�6�H�׸Vn�H��>���/ܴ��H*-퓘�!�<ҋ;�ds��8��<�����Z�V%�m��瘐,�n�.:Bl�)ѻ�<qML�q�����f�r��(�o'�U�$[z�!@8]μ��g���t��I�o�\���h�w Q	�N9��َz�:@�w;�����|�|ɐg�:	aP�D'K���UY����5љG?�b��9���G]p�{�w��0�D���� �36�]L���3��ޖbFFLP�UL~��	^�#)�Z�kp��I�S�p@�O��<� /��mb2;�Z�ͮKI�4?j�8z!���v��˴���K��>��o�k)~_�^.a�Q.�:c����<��7!���p���0�<�//H:�5S�����Vu�ڋ�Q<�3�RdE�C���`�Q��c�2�96�Z�)�)�-����-��	j���Wo��%9/jØ�ѓ�r��E��ߍG�ޗr6E����gѾ�}cuAM^ʵۚ�G���f�.�A{�����\;�d����f�SŸ(�hs*��iB�N_���.��-�d���+���ɦ�aק���� J]��6H˔/`�n���G�vk��e��/Wx�#�N��k#�LN��r��n@�L]\��~"�ux��~�1�!T�hh���q�����VQ�Z/���;�b}K{�<;*.e���EB�����+q$f�@S~��omќ�I�``�ŋ
fs�ĳ���,v;n�(1�� �%��׺b(��H/Ў����yG�Z�P�ho�y���@1��3�Vs8Ƿ��S�56*�t�0�Zm)E���E9��ԛTϜDC��qn[�la��*��4[���X�8�>��P�p���Ѳ;���=BGJ�;��n:�d��6r�uي�|�KXwIE�bM@������l�x��홸#�[�4���S��'��Tcڧ�͊m<�����ڢp�l2�[����xG���Bw��E
�����^�-�рFd�j�ҙ^�D9!֫b�9�`y4�9�$���Hb�<�W;�P�`&�oЕ�N
{\�9U�D��'�_���F������h&��׽��EԎ9��If���G8:�!�M�m4ȀcQ�����A]�>u/t�0!jQY?[�{Y���6�px��'�
�ж��֋1Z���6L(����rn:s����%�b�Y��������k�d�W�������	A%_�g;4�Ę$��t>o��3�u�ݲJ3����B
���H�L��o��R��r<2����q�`�#gNa��׈�R�y��G����ǿ�G��R���"��ϑO[ٽ���U�}�|���N��U�>����
v)��Kּ�0�_=�_�B��6Qb�f��ߕ��%	�ʌlU���5�R����ڗ��(���]�Kv�O!�-1+��p�O��TW���(|�SOxc�)��%|M2���(��o y����o���~��{r��Ȕ���J�W}���w$�՛>:$p�p>gm�cc�c-�+o�[<�}-��c�%��!H+�?��-���J0Ҙ:�zaZ�պ_kˁQ	��d�$�Rm�"y�ؐ�₯�'_�2�ey��R�����ҬWZ���7�L��h!g���g���HB��З�_���r�-"w��ӃE1G��^���x��A�I�{�4k]�^/x7�f�X"���c�,�_;��צN��k���u�����fgz�\]�G�7l�P�`>�{���s`F���UW��D�5��}D�S�X��6��Eۻ]�L��&����ƺK�[���t�=�gƾ)h&-��k���K?"�!1�mUg�W;;�2������ |V�T�N���#ȩ�ib��f�D�O�L��%Q����͆�(/�-��4@JDȽ ��n�h��kh�>,)��/gmA-j�p���g�>��c~݈E����p�65���� m�K$b74�԰���A�*u�ә��um�w���+��O�}�աl�J���t��e$_L����;}�'3��)�.���ߊz�J���q|�l��\F	c��#��f��0<G����7
�%�Tv�@�>QXwc��բۡe��S�Ӏ�Ά��!�v�C��c� �F�hB���-���a	��b n�r���F�b�w�>���i��0���kj��������]zV�h7O7�1�+�0V(� ��?�	�S৬�@cg}L��x=<�7@uE�+���E�ʤN�{���dv�Q&N���!�K� ��#]h�5i���bo��]����Or��t����1'f�iJ]��,
��p�G��XH�E��?J(�Fݣ-�����$z{UGxv��ɉX���8�� ����镼�����o�AN�W0���#U�>��LN}��
Hq��uX�����40 �@�!	^�B�j�}j^�n�G�G-c�O*�l~��x�{���,�9���B�{�x�_���on$1nk\9�E&��`lҥ.��ql�F�K_�n�̞ ��HaT��������&ƕ�C��KJ��p@:m�:��\���l+N�P:<w���:�$�Z
~ߛQ��Ҝw���}�"�+��@���4�O�xD;��%.B�I���BK���Aox�"1�r�:�"��\j�b}��X2ֺ�Lė7�yc�~�Xl�>j����{���}-��j���� �Į"�/��G�M_#C�yj�xl+2���]q��_�Ma�Nӄaz�߽�]��+�ֿ�a�쑚�l�
��i��L�@%�(f����x0BwG�q�g��C�9�z}n������#�V=i1O��K�Qc�u��,u:K�\�9���!\sBp�&�gb���yY͹Z,S��ߏ�~`�q�z.E4��u��<�6SC7�Y�Mс/Ӵ"�i�m�U�� ��9�׿-7ա�����}4(����H�o/����tc��3=r�f:�#,&�6�_���AҪE0M{{����aY@��ÄM�y-i��p����?��f4/S	"b���F�GUOԩf�NPs���
��@/ت9x�z,��+;c��m,{��[�Z���59���ȧ!�ڛI�:x/*�nHq@�9ɶ��* ?_�k1���z�)���)�����t�)1�	h� _n�w"�e�p�	1[\�>`lpuyJw��?"��~t�~/x�Ȯ�&�1�T�a8@�C�=��S4?��PD����^�"G�<� �=��S��^�7U;H�-1&���:���/��'���HڝgHB���<��3qrݚ�2��I(B�{mb∦�TR�"�������z���.ї�o�����X�>����2�����zx�#��R�ph�l�B���I}���#
N�O=/�q��t��5gˆ (��ǧ�"�����]���,E���Q�Y-��u>��'��2j�#f���ĵ;Pt��\��, R#���R�z�-N�Ndm��lq�������V��2�%X��.�b�����)�wr�=�q�*9�?��t�a	R��&"Gd{��`������Ce��$=0 �@��G����}�E���"��� ��Cq	�-+�i M�Y�9�R���H�''GE��]'!tF�0����}���D�Ɲh�},��v��������?�غr��/:!�0r1��2.t����Z��)��m�9����0��,�����ׯ�������c[�� ��u|W�t:wN����_ˎa��Lw6����&�Ƽ��H9Vo����6Z����ԦW~�uN�#����,y	��cA��{$�3�ʀ؄��Lb��Ø��h���ZM����A�6��Y����jvi�ߘ�NN=�Ґn��8M1��)S�2���С�ÔU�:��M17�>��$���O��&;5P���������u�x�_�c.�C�UR"�����-U<�*P[�����D'��Y���Ş��-��:!^(7���?��!^Y:��y�b/���Kk�����E~l�8~S��Vo�ԞZ����x����i�Yl�P�[Ȣ���I�g�Y2G�
���/�W=�3���%e�h��A�j>/Wan�s��k!d�޸��l�E��2=����}��^��
���l��?��u�(Ɔ�����B$sE�U%%�[��W���7�=��s�~]�X#�Qs������m3��$QD�k>��q��'ʹ�jW��Z�͙R搣���[�k|��bm�2�n��_�������\��d,�jn'_����
YE�[U�%������ʱuAd���F���X��n$��&��z#/Ø��2<�*��-��kZͬ�	JH�֡c�=2�9����]������uK�����7�S���J���ڋ=m� f�RVD�"j�e;-V�]�4��Wѭ�,A_��4��ĭ�,D���m�QNbc[�U:�x����u
��$\V���Xp��٦�x�<J�D�-��N}+~%�K����D��j�F-�'$=f�o�;��&ix�mGSM�q�m@�n����!��4�K45|w+��GUu���D�H�m�#[�x!� D:LDܭ�v*-)�w�`�U�$[|r�@bS{c�ڌ�,H��m_��&��W�5=���?c�s�i:�[���T婟ulXiI=�D�m]�@��͎�^����ɗK��k�X��vԾ��r堜�`�5�ػ�ȺCHm	�M��P��)R�ۮ+%�v�l��p1��5���Ţ�fA�~��ÜӆUME#܍���*�OʒP��9P��#�k�ߧ�[��KK�s��w<�/��⒐>�+���V��|vϺ��)w�9�J��5-?p�i�B�g>˷d`�d\V�T���~T�[d�T��&�:��?;��|>+w�8�6O��F�"1��r�i��5�uA�6[2�hj�&�u=����5@��~ ) ����R��w�O�MS��M��v1���r]�����d�)&����"��UOW�{bY#5�\�x]~va�}{<�S�Q�k���e�jM�-��7�n.`ws��j	����뿌��=��@f�=�b�>V�SP42z�%m�,݆�@�.,���R&�(y�^n`M���֙2�*��w���� )'�9���W�%�LQj����c���%%I�u'm<���q�$m9���a&V;v]���J0�17w@zD?��]Y�9AjB���o^�^򣠸Z��4�ˬBBR�� �i��$E9O��;�8O�~�9���I�a1]�&��*wY ����"�����P�)%�����t��#ߧ�nH��2���E�KM�N?� �K���񽾛��w�$L%��mi�X�a�b�?E-WM�T;��ʇ�O�)G,����Xv�w��Hb-�n��%u9�B=�f"��\�
���