��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1�i8��CZ�0@���}���r�$5M��{I���?��̱�����q���	�M�U�&g���@��,&��&~�/��G�*���s���*c��1�+��_W���]�����]�m��U�ˎ��H��'<7r�č<�E� �����������H�ǜ��ܼ����W:��4�>$��|��HG���o���fр�%��C�y�T�O���u`��3ۢw.��K#�x�s{+�u��w��m�t�ҩt�&W5#��L��@�̃=��T;d�*���A����?�繃Fl�	r��!�<K�c��%�7����,gOT�=8��;�Zkx�$K�}�}�<G�M�Nqv<q� �F{ed=;p�/I'���`48=���%b*��1��'��s)��:&)�m����Ib�tȜ�"��eg�zN�Օ�Hjފ��5�w��6CZf؉�R%���HL�z@X˰�l/�Lw������BAv<���`@ah����>�ֶ�Ck�r�ho8��$0:�D�KWԙ�} |0Da�	��G��~�u}�(�7�����R�`x����x�Gh���J	ct��wsQ�e(�ԓ3:D)$7?�p����"�S����y*fް=��y�����_[h�ﲨU�;���ov�~'~3_�H���"�T�������!8�"d�E�E��Đ܏���\O�������s/���o�3w3�܇E4<��0^4��ʺ�^F�Jj��!gmm�
}A������	g��`>���ZC�t"x��Bp<?x�V�� �z��*��G潖��c�Wrhd��:��G����p�#����M�3�X�$zc��4�F�.��g�]T��4�Ǌ ���àP�G�.T��r���7I0�ߛ�L�F����p+f?�5쁌���Y�deKD�����}�@A~χ��p���V0)���v׻���^/m|�����\�����&��z���ǯk�&t�"�Lѯ���aT?����ub|�5�<�,��.n�
�Zx�j�2�u��m3�l�0Ah½q���V%���q)���}�&i�}XyU��������)7V���>���MQ�ļ2l6���uȥ<4v��H���`��%J����:���4~NPR�G�n,9SP���^�1��3X���)l��|�L�(Y��%��s������n�\"?��H�+r:r5Q:	�?)�쪼�w�?�x�����&�(����BJ%�����֮��	��>�Z	M6��PaI�\��qe�=�"�K��h6���L�������k\R_{	)ܨꆮR�洹

O;	�q�s����P���@B����ԃN�Hd�<{]	��P��%NNhه��g�{�9�I��QJ��"��j���W�<��3蓼g�
dv��"G��,J}�ads{t���f]����/�. ��  N"^:�_uW�*�q��\ܘϦ�&:w�XmB���$���uI�H��G.���ا=L��%�8���4�9�c�Q��;�hB����-_nU�����[�;�	kL�ru-���Q�T�b�*Dq�}h��ʬ����#h>C<�����,2��a���x��A�)������=�z�'\�f�`����*܀��]NM��� ��j�Hk�{v$�&��w��1��F���⴦��0��8�N�����Dep�����+_�LQC�2�`u���_5��鷱I�Tw�!l�R�tn�B���A:�����Y%�r1�ڿ�o�"���16�۴ߴtR"x�T�p�H!�nN�W�/�Cf�2˶�)�R�]�Υa���f�u�	����Q�l��Cn���Kmԣs=T�P�z���i���L,9}�{7^s�di����N��<!9�$;g�p��)y�f��c	�&�47u~b��qs�0EqFL跡udUO��鳭z᳇�G��%3t��.�����/b=�̃ˇDI���%/��������l�u����2��/�p/�.���h��d2`Q���s{�1r�Ͱ�iJ����"y��ܺJ��:�0o�C"�g">ϩg��i'�f�G그�$���L�y3���	c��f�/����M5����[�L�&�,���vϯuPz�:��[���3Y�FP��ݒ}�rS�]��S�.y*YY"A����ː��D�bF�T��*�6�^�V�Y(s��|y�:rq3g�!�t��P��{�-���%�	B.�گvT����TK�����3�ɤ�s�����疢Q������������5y����Z�-E��\I�G���hJB�+���=<ܠ��O�n�