��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��]'��֍�0��3���F{y�L��u%c$˺�ÛIW&��h�,ĭPj�ԌF|�R�폽E_�?eJ���ק���Y��fΟ����1)��cGV��#�:y$��a������9.����{s&���f��)أ�*�l�z����ٹk�aNd�u��w_���H�d6��#�̯G�lfԧ3�W��<���*ę9����Ψ�WK�� �v-���=���yjMބ��{���Ow�2SY�<)&�#�.��.t�#�NZ��>xC����	�Ç"@ˋ9�����P��#��ۏ�nZ���WILz�?����|��0z_�=�ߒ�`|�Ee����a����f�ʓI��;0��I>��Mz��*ͳ�̓S�}�>Eσf8b�M��u�,��:�#�]��}��k�З ���FE��7��i�L0��[0O���==�ģ��c�3�X�c�	��$�ȐG���\�I>�C,!�������{��Y�S5�������	'�U�.�4����P��ЊT)�/��Y-��c^�����I�`�p�Lfn�����
�}j�3m�e�}n�@��|=�r�gPg:��2:�ϑ[��~� -@]:�Mߗ�olQ�WD
�V`����?�U�'��3�E�.�H&m���2�uN�һ��8鹜Z	���f}�-�:�v���Z�4uR� �� C#���[M�Ko�;aV:����-FKP��u�ݥ�)iXB]��Yj��|��`�%�[{�3U3x��XP1�k��ͣ�I���Ov�᳿U���4��^�(�ʀm��P?ۆ8<�<$�Ȳ[L����S�[��m���P��e�WS~n��Q�؆��y�<�Ѹ�
�Xw4�Dm��ggiS�Jg��sQ{���[��uR��u
=�K�C:�lU��/?A�da��%�Χ26Ϗ�+�v����H
�j���
�'ͷK�K�,����)@TSl� .�Dl����{hE9��zM�`M�-�6�����IYH!�o0[*cD��Op�wC7(q��1p<#�w:�I��M����a���1����o� f��PD��B��>���b�.���9��Rt��QQ�dX>�#"j��M7"b��͊8�!s��%0��%��~W��o�t�c�̳J�<N����p�rw����]�X|�)���u�=�D3MU��F����[{D3������5�CѠ��8�f+�����\�]�µe�|�FMk��;�#o�^�"�|ڵ$����n[-���2�.����.�@���v���N���?��G	�SM�޴��q1�i��0H�Zz�7g�OϴCm�~�#�~fx�zg,�V��<%\�� ����n�]��J�=�xvp�m	��|��h^[��W�/eUŰK�2pF�7"�I�(���TY���n���� ��r��Y"!>!��_<�ԋb>F�"�-#/�o�N���c%�8aoF�QEq��Xy���yW�tyeo8�1�����G#�����.������Anޘ,t���O�A/��!��~���`����%��	��)�xS��@N�u1IS/S�z�W!}���A��Ǜ���l�d}{V�s��S�/�tPd5nH�H���VHu3T�;sՃ�f�B� ���$O����|F�M5��G�>xq;4o�BOh�#�ߢ��䂌��F��!f��a���	 O� ��o"�Q���d��'���rά�-�~@!�z�!���|����E=�Ƈ'��~(-���١X��P����^��`��%��6�y� j�������}Q�����wP�C�%�?5߳�U30��	�Ǣ0Q��Br��H�����dp������,��Q�7�)��l�E�D�'ʓ�$X���`��b�����(y��c�.�-�S~B��L`�@��i����ԉ,o$y��R5���o���6WڿV>m%��3�d��m���wپ��:��2-D������[�/Q\O�n�Y��85"#��J:��Si��K)�C��)69�8���^�'B��~CsJ�z��od�Q�ŀ�;I��DzP+@C�����sL��R��t4�Oƻ�[Uvѩ����E+к6�����g��@�Vn��Sf��9,華�W T|�s=�'HU�6&��Cl��U]�����J���	�Ȅ.�Ykܡ��u��}�#��(��Ym�e�M�%��#M�����հ_��~�io���H�.(τ�gPVi�Dh1iԌ��$q�� �J���f���5��῭-�����{:'���5�:ұ�����R_��-�V�Z��K6��9B���k+����!����|�K_���77�n1&��I��ڇH�q�}|��`=��V�v?��x"@�jҟ�����$\�,��dy;G(Lmq��v8CŚK�YD�XN����KSc1�i��z^kl������5#Y�qK�Хe���|��W��x�Z�MP�f+��ߨ5Q쭿�&]��;EKr�-7�JW9(�U.��=C�7�҉��®�ghR�?��}�0Q�<OG�z�y� `�|7LDk"�(��rThtU�
�9V�G��$��l�����%Z)ɚI�hgY�k���*㤭��� ����d���lw�'���=/�d��DP���	���okjۚ��*�Ͻ@�r��ߠZ���1�0�1��~�>_~�_�Ý�����ʣ/O@Jσ�ǒ����ZE��+19�#d�;=q�L�y���g���K��+坋�n���tUfc����ϯW��o�\�*I�Q'�
g%/��N�]����ϖ��A�G>?<�	,p��һ�.fgr.��J�h��R��1��K��㓬��e};�[g�+��9I&�8+4�$/8�"����~0�&Q�R �n�0B�ƺT�[B�]>�Pŗ��7r>�'�$�R/�Q`�(����j�K�Hz�E,�9��������t}�:u�tδ��_CW5�w�7�`s?Nt )[�-����@�.J�2����}�O�ݐh]���q�E���s?Ɋ6��p,�n ��KB����DY��=�5s]�"?���y����C�N[��,h."ܿt����8�Ƶ��MF`*Q���ħ�G,@���/z=cI�҅��j��粦�Е���wz�"���E��:��HU+���J+�4�B-%�X��:ֆ��	�L�2(��L�GF�H���,��{�SľX$��r6����-N!}���}�K�%u��N��7Ѹ��m��f�H(o���&S2Z���}�=e�M�F�'�3�m��f���2�aZ�T0鿩R�^�p���n"�&��������d-.&�ï/8?c�q9	��������?����V<5W𲞴W���U[�b��-�ob��|E�W@���h2�[�5@��1�'~�~7|�"��l�� T6h(�� ��M[����>�H�QB�Pr�u#����v��Ă����l'Aܱ,�-֎z|(�&���_	A���'b����{��m߽w������}ծ�H�Eeĭ�j��1Y�;���ǹ#sʹ`�ԴU�D�$�����_����'-�������A���Q���ǙbO�}��-��r��͆t�C�^���?�{�	�ΩŶ� U�����R��=�$�!���/ �\\?f�/�0}�>}fDf7C����ϼ�1=o�y�&Չ	��*k.���%)�;=-��>��@'�������R?���x���zd�%�b:���-"�7�K�_�M�k��m�Z�!��-�*5�%��M�d�i��T^\�>�N}�����/�~�!MBG�Z��#`j�贚���I2Z�����"r��&�<�}�T���w*ҭ<[�6o�x���@�A®T�65��0�Ka�x���F!�F�$��ˉ�V�4�k��Skr�����ۤE���fPf��|h�nyN�[�2��2(�dޖ�2�Ϸ��jcQuA�g���#N.��cF��%M���ӫ�`�R86Y��:�S�c�˷[r�Ne"�2!uіC�{v9��?����L���[�e��8x��?�^�H��_k��y^� ·/�c�y���(���&7��C�po~!� ���*�sJ����r��c����'#�!)�zaOE!��zn��7���P�e�6���o��1�;s-�#"G�`�H"~2�
W�C������u\�X�N�H!}�@��Sp�o������M#��%s-�BF��@����Ri�|J�#A���S�-Z�Y&�$b�6���7-��w(�*� �J�����f�Jry<{��M~�@�{রWj�;%H�i�}Ƨ��������?<U�W�!B0�t�L`'&�|y:��4�F�"���SRQ��3�oRw� �S�����bJ�x~��oG-p�������� ��*��8Թp��������5L�]������z�>%#��r�h���Θ�T2�1�̍Ѐ4��؂!Z�kϓ.ı�Fx�ߕ6X���k���0X�5w��%?E8�O:��z5;���؏���
������qAB,����T��Ȼ3�;��ُK�l#���Ƴn�;|}�-CXU�A�M���*���OVu�;��ߋ;h����A:���'��D�Q��]�"9���&gT�;5��֦��M�'��V���"��N_a�l�+����BY
9n��&V������E�\@ Sg��L�W��[X@�ZT��Ӵ O+訙qb���P<���">���� �SDm�
z�t��8�Ԃ��.���W�W$�٪0F����g�2�>4��Л5l �$�0QS���h��_��m�P��ڗ�蟊�7��Ց�n6Q�%�F�䖧 �8gs�o�Gna����D���>��]s$O��� B�6�!��[�_܄g�qb5��L��n¾����<��RuG�]�Ә��O|��s�Z��o&4��� H�YV�V�>:��:���֌o?%
��#}I����Wh(��!	S��="�n��V�n=J��.�2=�� "��P�{c~Vw��ν���N�?s����p7 ���J]>�$/�:��VrN�9��&A���f^[S����ͼ�=���#H�:
��^5�?~�rX��'x���{����z"Lc]e�%�%��b [��t�I�&�w�
q�Fz�N��˷N��ca��, �O��8
�3t()H��(7�E�&�! >i4����2�����Dpi�}A!���-�P`5�A�k ����<�%�d٪v�Xʘ�<[��Ա����3OF*/�]Lyx4���n|�TE>��%����Ag�}����~�G���h�
���@h����6M��9�yF�%X8e�^x�F�m`�F���lK�'��'�`�)�#�*G���WCv�Us]�u����p?8���AY���D��"�o����&һut���a;��!(哳yb��y��]�e}nD �6�7�ֹ�%܈�uh�e�t�:�����I�t���5�}�WR��Z>
� IM���]#:`�"����U��l[`����[�n�`#S���\���xB`��#�UtE�
�&7�bT;�@�=�;/g�]o�`��>�p� h�d���߷{����5`=P�R��%oF�!��O��id ;�(���~����-���1B@;���:�M�&���E� ��� �wY�" ��H���u�$��U/(Sհ�qt�e]��Z��z�����ݔ!�j:y5�qA����U�6�P�0nO�z3��Q�(3��\
؀��y�6i�+�E�ta��вҖR�wtM��<X�h���X���wIInN\�_a�儬��>���A�ӄ�_2��B^A���U��a����Fw
S��  -�����,lrq�03��D�3ș�zjr�o�9z��e��Y��R�K���P���⭮2�a�^b��^���¤n�"�a�ּ�#<���@�l�܎�j��I����7B�ڐ�?]�"T~s���NK,�P��p!s���i{A���s�����B�Ҳ<qa+kW&V����Ē�er�;ZS: ��+I�\k}9j�]��K�ug�[7��Q`���'�tL7���I��	��+2Ώ��jHX���_��}u���$�/p^�!����Y>�fc �����m�����&ɛꬺ�9�������<||:��<��?�&��jqJ��=���!�[��㚓&�Y
)\"�t��� ���%�v�eR��" Y���dAwA~W�#�l���Y�r�T�5�Q
���JM��Άm�[�ٱjzkzJwu�q�R^��jx����؊ �`^�$�h�;k;��$�FB�H���W��1hd���&�j��V�;���MϚ	RV1"�d]F��k�֪X`y��R茤��Gy�%�p�bR鏃�{t��f*���h�/yN�6���Nq'[g���:e�^�(�D՜KxS
s���ƒ�}�����S��(���'����=�5�8փs�(�Gz������V������yȈܼn��ՖDEKW�����Ix4���(�5m�7e�*��0��o���B�a�n<���#~M���N��?�+~��r�M������N�P暤�BR�r�����6��ߖ��W3�7'äc��\�:1��;;��Y$e2n�N	�q��Tg�x�#N�4^u�
��a��%ILiG�Qsp^�\���\��M��w<ß��k�F�1w(����NfS��;�x���9�t��V}E �K���#Qį=%
IT�	��Ͱ�/�1�����B�d-�0�D��Î���-r#B�yB�w�e�lS�Nk�16+����4�]x�ptuK8����vc��*���һ���T�t�Ʀ��Ɍ%�b�J�V�w:�nM�=���S�zeD�����7�y�1���7hF�q	����.
2�{t@]��{����!CN�<S��1����F����rC�Ͷ���d�2��Dnv ����՛��{���Yų4	��E*��@���(����Տ&���t�I�fN�����E�ϴ���hr:n���8�Ք9A0d���x���)Y{qSB-3�)����+��D���XK.]: ��4n5LL��lHv�{��WD��H�5F�dwV��PY��yK�t-�C��o���w�2Gr|�ʋ�X@H�Y/I��V�<#,�[�����0��q9���L��_�-�z|1u	7 -�:�n���!�v����Ț?�U��~3C�~7�`�au�9K�f�2q�8*��{��_�~������s�>���{���!���*Ӫ)15�b���������:B���1���@FK"��JA3������`��sk<��.|;,�C0��|�/Ȗ������q
CD�
Զ�=�p�G@aΉ�
��c���qL�kOnP%������7苘���pG��>A��c���Ek��Z�Jl�J���ݳ������=�b�06,5�8;�F���_��i�8�zU��OB���?�������
�\(,�3�W�H���L۵�c���� ��߹����27X'
���Au��u���t@�a犜���-Y	�����֨��yt�0b./v!@^��!��'��A�wB�ߺ;F�(�S�=V�rZgּ
���LS�aȽ��h�E�[4@�XGI߯\�����KR� 쳢S$�o�	�] ׏���'�$c�^~KN�Q��w�&�PT��G��n2*�-V���R�tu�������M��%%y+ܮЊ�u��
��~IŖ��������=��bF �V߁���K�VX��Nw�)�ۓ����2v=�1Z\K���5�8C�cў
�u'�X��;�U�z��@�dƬ�Gύ]-+���}H���Kv(��� ��ݪ�o�d������� ��.5�#f�	���](���:��!�p�n��f��VI��ǡO��)>���X�0�X���Eb�l��m�8�?������b��9�[]�Bo7�����/J	�C!�k���ª5�{��DMս�� 'ӫj�ihXN�^����8������f�Q�@���� b��`L�ǉR�tp����e��01��:&OZἲ�'��A(N/>��.�R���K�UX߽�37��^��+I�_2�;�y��*��O�@�Vj]�C��8(6�e�2�۪��t�a���Ex:��P8��A[�j����Č:�Niuwc�w��r��"Z����9�3�0�b���&5��~��5E%�Ws�6�̓f�`�B�}�C�7,h�4��_=��R�������4C��=I��%q�E�^��"��fvؓ��e5�z���p�"m�`�rD{�ce:�	zҙM��<m�ꛨ$+�r�#:��<�4�KH_OS��=�D���{Q㍑�mELJ�<�ъ��{��3�~���Z�BQ�'y��F����(��W���>�S�����\� ��4���5�zo�u����]ABV�0��V���x�ۅ�rQ�AV�M+-����@�i�1�ƙow���Ή�*=��\��h�q����nF�����3p�-�'ok]P3�>�P-�7��G��U���,f��#wܱBw�ww�,��e�(�A��n��N�T~K쀸�K
ޓw��1�&.9�p
f����Q�D����AVl��5�9
���A����=��P�!�P5˴�|}"l)~�q��يwοֆ۳��k
7�(�J��4u�V,m�<�>�#{����H�������Ze�<�Ess�O��P5�ۓh�yv*���+�)�F��.<���9E����,�䟃չ,��I�-����w��2�D��)_�(��]Q�)��������m��9M'\uf��Ԑl���撬1��PLB��)hKuc��)�О��t�6�`B�J��w,Ǻ4�镇� 2A�&�4���܅'�[�zI�F멲�l��Wb�YB�U0�I����?ߋ���[���l������7�$$�f#�E�-;|c��R���2[=Ҫu��2G�B}`�������g���oWr`�M�`̶ 9h+-�͎��j�5F�k�"�!/��l+ӽ�1��J6��U�)R��tҔQ�\���/���x�@�5���Ou��nT�� �P���C�x�N���Rve*A��^�B_[Ǜ�crd&n�s��g��Wx����=�A�=�����%p�!$��H�mm��A�7'��3vJ$u*ϒݣ(�$�f!��8h��=V'_���a1c�Bt^|�����/G_+�~��M���gUK��Z�V,\�"��P�vm51�l��g�C
�������Z��#W�Z<o�Y����A�>6?O�� �F��?Zd���߬.K�Ld�oɈC�F�ʠ� z]�*~{@�/7����bdU_,=���%�aC�:� ���[�>���~�FA�xA���u�V��_?��
�3ՍI{�i!�8�(�uT���n������K.x%B�w�<�������6���\l�
�
l>�R	�P�>͢����q���Pf�Kb!�.���Ɇb�z]�^������br�B�	�|1Y��U�M�~��r��$3$���јl���
6�㞇��'{���z��5�S����!��r��Ӹ���0�Q�O���ݢ;��%�qc�60H$[�l��D8e���S��p����o)+�ȐB�/YT->�ׅ빠��1K+>+�sՐ_��h�h�2w�Y>��_����D���ށ��Hﳍ��j �<�$���G�g���%#�=��~tZzj������+͒+��`�5D:.Q�	=�zN4�I���#�q�	�$����"Gai��Ce
?�
�n!_��59�6 ,̯?o�4�r�훾0�͡a{9�uJ�|f��R��B��Y �I2�&B@ע�d	,)[�e�2J���8���v q5���LЁ���"_bo�,�i�X}�8b�O��-m'm�d���i�1��4�k�w�U�f�����TmJj�T����1�Xu��V}��
s�xߌw�Za�,�c�J���^ޗ�����7�AQ�w�F�p.ɖ*��q�8`�ߎ;����i��#"F�o9����տ6�㕖	ݜ#ǖ�� ��ڐoO�r'��D���^�OMi��ʺ�U}�� ���
VrԻ �1�3Kg91��O~�j�L^�
���IZ>���9-vF�Ęd%��(2��H[���*�zpݛN�"���.�d]Q�[ԛ<J!\f��9A@}G��>��g�j;}ʻ�ۏI;~���^
w��2��QOhݩ1uwDY���eZ}4����ml�)H�֑���3�0�YG�s| .��ɠ8�t�Y�m#�8��9��>Gː���+S�|Ў���_�8�F.A[I3��-�~(�+,���X�r���R�3�h�ǃu��KQQ$\�W�[E�g"���f�/��ӨDD�a0,�<U$��'L��Ӹ\��2Z/y� C�/�iuCZp��]��#w�x2�W}�e߲�F����K���� uH��P���Lc°r����m[�#���~��E+���N�C ,�	V�/c�p���⢉E~d�E���d�?��� ��.7�/��L�Z���'[��YߨN���/ţ���^ƒl��
Ş�6��(��X���C��P�GZf'�*�b���èR�2�)|�IӯK�>�L`��=M��0�,�/x���r�*�a�׷�们�Q�����2��?�Q�S�����\ښ��lc�K3StH�,�g`��a��}X]|�^U�%�y���z2���[L�a��@xY�K����qE�Ώ��DF�8��L0�C�0KZ?
%���)�X7�ͬ�\��FL�Z�8�r�)e�g��.�˜�Hӷ����nuJڙ�.��H����P�"�T�]d��Z����]��!}�r�o��8}������_�V�+�����4����V��{BQ[�&1�336E��b��6:�q�y�Jhjm�����w6�.w�|�r�y��.9��[M,��NO½MϮ)�z�ve�����v Gc����3_��J�[]oQba���`JYTb��gn5ߤ�Z�j�$>?��n�
CbhG�6�8�g��t}���5VW�؏��5�"��+b^	�D���c�d�b65
E
:��/P.H�&�V#Fѹ�A���I�g�j6�Y�|�y���jJoW�{��`�nY˵E����{2Aہ���Ï4C1_Ew�z1~�s���@)���͉{�����a�қ9���yJ�JzL��w�t]v(~g7����)9���"|ꍦ��ހ/�kѳ#M��u�*��VM,`�/�nr�����{�=^�h����(�y�¨�g8��f4�̆����{�>e�^��KK²W�W��O>۠������zuN�F�5:�2��oW��]�-d����g^r]1/%�̡�'�}~�r��%f3-y�Ͽ- H��IE�3�-�<"Y�z�1U6�D��a�DX`\MZD�*�G��8���̭Ϟ�+�����P}��h��w}�c����˥nа'��TT�S��+-H8���	�K�$<�nm�ڄmo=���?��b��}�~I�nt��-�Q1�?3mv�����t��EmJ�ڐՏ�PJ�xh�Ч�^d��i^��-�������gkӝŬ�'� 2)�fj�i!��s��:�(�"��:�)%��4&�0�Aa�r~/ �4�y=(�rO쨯�9�˽k�B;�9�8D��M�.ͺv"�_6��3��MX|�8�]�M�}v����ڀ��H��I�b`�\�l����p~���%�~�LI~�a;+(�X�w����<�W�~�+z��оs	��E�Y��a%sp)�h�޸dd�o�+q=`��V��I:��TVp4:��Z���n�ڭX5y�@Ы�����"Xf|5I9�t�1m���iC:҈>�K- �݈6Ϩ�<$~Gj·�h��!՞��u/�@������h�ﴲ��C`29�Q1𸡗�`��9	�Wd��_�zu�;�����l�I�-�F���p���{+��pC�.�f�`���̀-��4�Z�\�����Һ}���z�\�S�.lM�?
%��v���ۨU��z�b�{nL��$�7�CR���(�`��_Jj�?��L,��&W G��D jώ7�[,t�%�äO�W7saI�c����mRU�yE� +���L�����͟H����w��cw�t��։CFX�&��d� ���,/92��*�M4_Ӑ����%A�F�خ�o�"�QL?H��>�����Aa���.��61:h?�݊�����_���52d�\u���<���@�	M��5��C�;��T�IӼjy�Il�Q�����e��:L������xDq5�0	��Ǿ+�/�M���y̴�₹u�A��O�����J-�k�!/=�����'�<��AL��w����c��9*׫m�Z뾄�~��iI��^tb��N��ax�8�9V�bĔ,�A�w���)��'�m!)��<-ʿ!fi�a�#��>�Y�|$3���A�*��Ȃ�����&�S+DD�AXBV�vd�,�<,��!-z~�4j<�Tl��?��$�	ȡ��ݹ���Յ�1r�ab�Ѭ�?d�MR�3��'���*Gך��6l���A'�Ar��D
� @o��y(&�׀�h��-�f8�i�����WWBdU=�8E([�c�Q�a;��Ι�c̹��.�ꯜa�A�=+O�_����v��42y�D�,\�l~�v�6EC�/\����n��=�JV��u�l�r5�Ĺ�f=mIƐ�/.B���\�d���.7��j�U*���j����:F0F�>X�k=�@�lh�m��wWM[�6���'�	�Ք>i�gCPa&��4.���}7n�R4^Y��N�|}�1���R���n�t?*aR�Ǐ4ȕ)��R0r�@�7;�����y�K �(���_����t�g���cF���`�W�|'��,H3��w����Ҵ,g%�q�)O��*�����_b,	.#7	b��f��f��=��k^��İ3f�E\9�G[Mӭf:�6â4.|!)��τL�Qҹ�g�����n���+���&��\������r��2͙��tԪ�س�Qwn�sE�1xH���[P\�3'�x�K6����Ɨ��ގ�����d�)u�Z�6�E��wB�u������=��;W�tU���0ד��Ί��#����EK�x����`���)��[Y>#9T������}��y��Mܳ�al ��;D�U�ow��A�03�l	�Έv� 	�yV&}%���O�R��>���J$G���۷"TBB^|��`	�e��E�����>�߷W�����,�����V��?ތ�]����4��م����nM\r��ԝ1����	)��˕f}?޻o�W(D���.a��g��l��M���Ji�H� �זň�[��W����K�E

��dW��~u^��0��P�R��B\�P�ʋ/0�-l�����}�5I�:��m�ֻr��;	�sSCw�Խ*�y�k��}���!�#?�;��ԉU��N%��R{�(�������#��'�ō����+R"x`l_QG˒X��k1ψ.�!Q���� �)����G��p=X�C<f���(fG�κ���8 �q̴��R{�7q'2�C+O���܁1�J��_�}M����z�\�v�J0ω$����8o\Wa^�jF�o��		\�Ӡ�1L�}�-� ��I٨�����_G�ͼ�4ʺ� �q�eӾ9�U�ehߝk�l8����ҝ�3'����mA?�%1�k��*-q����\6r⪃��{�1�+t�pHE� ��F��銼<���Y4��*|�����c�=� xx�h��&LȠ�>�#���oTa1�e9��	��<���rbT|�4�/�|��Zԅ���#;����_������6&t �)x����� 쓈T��/�/Ǒ0�����T]�4�v��,�Wo�Y�:>�5v����GϒP��[łz]��y��������$�h�R(2�CL*&����d�c�h�;2���?O� ��BǺ���.�Vt7��E"�1_v랅|���,/���҈���Ϊ�� $�F=�Y���}VG������)�_Y��̃��v姹�ANj|8��I��p{7��FNld��4��w�4���D��H��P�p��c*FYǉ�5z�{����5�Z�T�t�P���$R�]����6}��Η�E~x��$�]��M� ��@ ���q���5�H��/�,�Djy�?VUŀX�75�hn!J����6N�2QB��]]z3xb�D����;�
L�����G i�
�ͭk҃�v���Sx���m9w}�b����ak���@H:EG� �e���"������pR뒽3�4�{5:`U�SY��lt`b�ބWn-t@Ģ9�{򪁋�Y|�`7����Z=�{�����2�AA�=�BT~���K޴Ș|װS]BkP�۶	�4;����Y��Lj�&��ã�	�J/��T ���ÃB�i�\��v#�0�X����K0����az�cE�_���a'�B3jã���:̈́�h!r0���
>K_>�O.�L� >,)5F�Ρ{h
�f������u�٪��_h<��u�@�:!�cDa�����ސf������G���U���c��m�[�
���2	_�������D�;��0�sg2�5V��Xe�$�~`�!;��y���A��蟐W�c�ۑ��+�Pz7&�*N}N���A4�g���$G�� ��8Y�_�f�I��a�ܯ�$�/Šp��@\V����z�'�c�V�I1S-����ϸ���M�|���}�*� �D��@�hGf>�=zB<{�tYE���1���[�Oo`omY$�/�̄��@K�i�"��{+�;��D��"�::-v�dGK������J��gΚ^z'�V`�75���߰'@b%?Y�|M���)/�;�m2�B'	I7�p8�E9;�D��� 	�]v7 �:��B�5���rکٻP��Hv/y�5��y/���D
m���Π�k��O߅yV�s+��~(���|t����Sn-�&);��@}��	�WV�������㣭����o�/��r�E������H�C��h��>}j�wZ���a�:δ���ne3U���b�!�C����h�Jr-�����H9(�ʗ2	)1٧M8�5��F`��������������b�W�w�kl���;���6,���aL�tc@#��1j��v�-/�=�gt�1M�3K$[�N�sկv��?�j^Mz��D�
�"%`��ٴjk��bl=�64�p������/}=?�!��$}2�NW�b��Y��Y��0t�-)Vc&^�@���`خ	�`��}i��2�u�|�6?��R-=;����]�X��Y44�ޛ��j�Wm�
${7��"W��,U�,r��!7ʫW�q�~�oGp�\O�.���Y_�8n��������Rn�0+���*�:���Ʌ
���P��d��	[�zJ��D�o��?� � i&-6Չ��b	'ZO�<io@�O����y���8��el�L�錙'�Q� [$�P4㭢��oھ]z׭~5m-d���v�s�t���f����C.Rn�q� �����^!a���g��2凼uM�����r-%ۋ�S��\���@����ݏ�~
fOv�V.r�a�A���!mZ�JgY�k���%�1��Q�Da��M�;]r،��K�Ȍ'��0D^|���Q��%�ɡ�=�g�ɛ)9���R���ۻ62&dmD����C�&(��;�G�����e�f�=ۮw[��!t֎�g��+Rәg]NT�$[}��տ�)U<�^�J�y��*��4�g'�(Iյ$� ���z��6�M�>I`v��l�XF�����NFH,c8m�=��%nXV;���ԧGb_W�� ��[�F2�̧ٸN��?�g'�����e�Cp|k���5��u��z��#<����2e�w�����Dm�|���!	���,�=����C
�s���yOd��~�x�'rbҩ����L6�O%�;��i�ZxȞ��[�PƠ2
���ÃB}GB�;y�y&|�u�;6�`Eb��i,�Nԉ��ޘE���i���(bP�s�6��p�\F>����V�o�c��!H�@�+b����\�Sl�ڰ�HZ�yE�d$\�N��k(r�Q/���5��k�_"&2�P	α�2�K}߃�C��՞�W-D[j-:>R�E܃@b��������WN~#��9Hѳ��)?�t�%�@`a�&�^�HG�sZ��u! ��>ϽRl܍K ���!��Y�w�^��^��j<$�V$d1~�e�L +�P��DZ���)|���R�`ό�_����}����W7�� �v�a�R�0ꁳsD<r���9��j8%[	e�.��p����X��6G+8�E���&�]~H�%m��hf�0 �Q@��������_��F�[��
vW��oD+��5��3tH=��]���=�쮤d��%�1�V�|�D�$:^�h� SD�1���[�������g�,�	�f�[��O|E��ѧ.�œ��1�Җ�FE���M���.�K����j�|I����U|���ص7��Y��S_@��Y�N�#����s�^�'��ݼ�,�������>��d6�mP����#G�_�kD�p0K�C���i+s핬n%�L�c�&Z�D�ص�Z�#p�aS�d���q,����ĬT踑%��nf�馶�����m�rY�gA���~w�����+4�,��$*x
ct�'�2��s)f���H2�ݗs�t�
z��T�t�ڦ^��kibP��`Y���F!�ޡ�ܗ?��8�̲���V�#��&s�Q�R�ll����� G����6j�����	���x)�
���CdZv�������F�X�vzi�,^$P�B����4�%��{�D%[t�t�$���.�3.�t/
~r()vQ�����C7ڹ��O��W�>���w�{��:!p0�ڸN	�1��7�q��zy)�ët��ƋO �T�0O�47�f�LAw�R���/�M��&�V?�p��c���a,��b2�_��դ����}�>I9Τn-{���P�'j)��T��X0x�[��(]]'����$�j�\0⡜A [J�쫏`�������COz'Vݢ=���8��Wq�N`�X�}�����Q)�c��j2ʚKg�z���PS2#(��E�#���h���Kklc����x�v�`�a72yp�_�S(���+&��1�~T����a����y��wO �q��yL����p�og+��G4�N��Jm�A<���)���<�twR`�2�B�U�.���m�x�BR���p�4sp��"��n��=	�)r�|Z�|������PI�'�aCf1�+$��B�/���O��_�2����ӸI�&�Ӄ���~��}.Q,F�#$��ͣ�v�+q��0�~RO��x.��􁰊�ޡ������l
0������s�y> ��[58����������}�v��H��R��nw_MD��v�Ȗ�����La�ꣿ�&�m�hW^y�����ԣ��Z�x����B /�Hg��Xr�~��ǻ�
�0��(��[�q���օ��}e6��*��O���3�3kR�։�����%�s��V���"e�yw�Bp�}�20�)P�pA�)I���1��.�94���y�m�燰��Z�ڿ�e ot,���~���&�TDK�@��#���X]S+�a�IEor���a��2�G
��$ diQ���E��I!^F��Sݨ�i����U�(��>ɣ��dl���L��h5�f-d�g�0��б0DV,����<���UR�x(�Z��;	�I5v_�\/c��]�{`��V������鈉�#h=��o�C��0rE�ۙZ(8����J��'6	���_nΏӍ?���؃�J�%-��Ӏ�^�z1w����<P��zmA`��}Q��iﱾMI�e�N��e�O��C��i��	E�E�ߩ�)��Ch��]y9Ӣa�y���s����>��Bb�SSZ�.�&H2Uذv�Q����.�J�@h�Sb?3���+�I8�JF��R��Sg����<ǫ'ĉ��D���B���]3��
M�^�6x�ê��q�k~OT[ED����K���7��V��7f]����R[��0��Ѹ�KjL@�����%�r3s�ڴ�l2���f}��Iq(Rj��Y`;gb-����oK��B���;B3�Dʓ�>@x5v��a(!��$�� v�-��EGh+ꡬ��^�9$C/�*���%e'�ɺ�A�S�^J����葇E,��L�2|����Z�9�����n����D�k�*(�u�^,lR:���@ُ
οQ	D��MJí����6�	��GC#9^��.[.T�q� 5��]6�pd��q��eg�&DxE��䢋b�͋�H-���uؘrC���o�;ƹkzϱ�?PDq���R�\n���G�W�c��#j"˪�/��H{Tܳ;�R�k�]��F�y�̦(�?���z�G�6?�
�����(�{7����A�<���+L3VRi���Կax�����{1��wY�2d�LeRNesuȎ���o��+q�F�yުd I��oln�1p��OU7}�ZH���O#/\�5N)J�lo�]�+�an�baS?��꾺��d��n{�z����!T�R�d4��+�u���xU*�b8�o�&�^��81�~@NG�:�#8T�E1Lq�Ǿ5{���w���S�8M�"�p.�Y���@�i��g�1��*�N��L���E��� ,�v
�Y*<�S��y�����2CkI�e�b>��k 9�q�Quv �D�ς��Wy	Y�)CW�ʯ�[V�8)�A���5�/��L�;D{B=΢��y���n7|Gy�6�Ū�N76 d��<�N^7Ъ@&gt5��\g/�(��j����������֏�QOJ�T�Ȼ�畘�7 ݢO"�s��/[�r�rh"q��k�C(�s��&
�wc�&3���97�C7%?�������o̻C�&C�s���is}3�ӭKU��/S��t �B�0RI�'�D���(y�f�,Ɣ�{l9��;
J��^����>L])��Lq')��o�1�>���&h�v�S�S~7t�����i���=ӆWy�p�>%}-����ŏ�:�J�K�x�z�sHgk>oF"��d�Z
E�,�ݥB.���y뫅�+�0�B�(�͋�K��J����Oi���!�ݜ{Gy%���뚃M}zH��g���OV�Ov�S�N�7N���Mv�O�)��&M��Kj�-��������B<5S!%��u���蝂x��j����h|H��"_Y)�,F
C�� {6%�����<�E��pw��!(G�E��a�Z���kC�
��><i����7��.���n� ���yr��ZQ��2^�6w�����9�gg� #n����w��H�L�L�@�K�x��[�d���	���1�쓓<i�[��F=h�	�zm?UZ��t�׶�s\�V
���T�qu4�O7M�q`֊�[�VΠ5�#釔��aT�̨�_� a���	Vቿ��⌉��?˱�Z�M?	��d����^�.鉱>H}S�i⚏�gq��&�K���V�je���D��X\E%�gO�>4g�Gt_� ��1�}�dɀD�Zt��
^鐑�ԅ��[o39��ލ���U�y�G�gW�'�� r�S-쳜g�\y\����/=]�Qʧ���$�}s�1)U�̉LJ���aS؁�7����c5��sD�S@5���N+5#����x�w��4G/R��d�g��87�
j�O����Ԡ�6�2���@��˻^���L��dLs\� 9��~�*6�X=�6˵�_  B�Ցן�]�RH��l�pb�����m(hq��nc2%�7D?�5�&Ü�������H��c�kb�o[4�n+���#e��y��K��,-)H}�3�#��0w�2�����bcm��8�CɆ�-"�K�q��uz��8��ŀT�R�{���QB> vDB�A	(R�M�}�B�(�kfr�pL0'��i��)��?Ay�����:�?��N{p�S��GF��sͰk���j����y�+ʾ/ ���&�OKB����V~m`���7뇇��PL�$(rH81���R͕���Ѳ]�N������Kl���iW�a��/��Ll@KV�����|Cu?gҷq9;T�K���c�ސ(�b��I� ��e�ܖ�9��7	h���*O|6;-�{���NB	դ+Q��+~qs�Jv�Qu���@���̼U$i���FI9�c�%Tx�s4N&��d;���� ������t���S�A�3qf�JR�і8���X(y#��D��!�I��|�^�N��jÄD: �	�M�V��{+iR�w� mQ��i&Ix�����5m;��%�f )Z.�˚5�8�_�b�&j֒�\3Y����������enx�ʷ�R�ֆ�����ߒ�~�����x��w��>)W�T���Ee�I�ZZ�fH1�!,Y��P\�h������e�,m)�NT�9bmͪJ��Fٍ*N/ݯ��ԑ���W��hɨ�1��!�#�),}ˍ��M#�}�Er96tg{��V�34�p+.D`-�C-���HYv�ђ�d���������Wjw���!����~�[�;WT8f�8����c�q@0�u�sw"��֨Y#�7j����N�B!՜���\=�8�h��L�Zk�0��R0��g�_��I�u���Ĕ��zK��C�o�Q�>i�^w�4FҀ����ǯ�1��2W䦞S=�Ŋ���^��xz{���ީ�c�w�r�rƘ�g0����N=����q:v�)H0�:����u�XN�$�/i~6i�Q/�4����@��A���ܪ��k�k�K�y#�4�@Ҽ�������z���	��^���q/:���F��A~q짒�^����&`&u�^���������C�������|.2n($�hդG��Jf3I>���C�� -#�b(��S*�_l�O@l�<x^l�0A���I*���8X���F��{�$�K��4���Z*�a�2~�i��km�5�� ���t�L�=�fR�K�������oD��_�[��--���ڌh�Hk0�_����Q�p��Z�[����.��I�p��Ai� �m�6�'�k���¼�B.��<�d�y��ل�d#�fN�����9zڰQ����%��Z�:����ҭp{^^gPT���m��f������8巹���z$�#=/"&R#��V���F��S�7�X�@�,�S�L������s��3��ex�bJ�s�,)��6$��I}���O��`�����H�-�M-!�&k��j��Bx}ʞU#ѣHv��)�Qړ2k-�X�g$��%]���M�G���Whr�;�5��Ld�rA��KIT�t�p@�ql��ON�O���!]��#�J�c�*z,�󢈓\b~u؈��!��6N�,�ٴ���o���m�>N�N�m��2%�T�h_tx�x��8�Ԉ(B}��������-� �mFr0k�m~�;�b�h�b&���c�:��]e���#B�q8���c"'P5�n���]�Թm\2�6�^\����A���.�wZr����8/� K���R����=�;j{9�(�������mMm�@=�����R%=��a�����x�
��f�/�u
���S��}�����͝z��)vH޳���o��|n�Ȟڈ������jB'x_@�ӹCl���h��4�{�c_
	�i0R��΋��[��=�x��_t8a���k��
�Z�O�C�	]����JF�Z��'��V�.��Y�q����l��?�c'���~�,��Y뙟2u������BKDɏ.�'���o�-�������4�3Ѹ���?<�݃�\�&󸵤�:�3'��>R��c�/�Y���J�^_�W:�����B!���ޓ�`L��E�v��NmK?4H�����O`��1U���q�'kz�)lg+:߼�^UqЧ,/G��튃L<_�2XMM�5���1�nG`I7o;T:21�UF�LC��d�Qǡ��x�Wݛt#����%9������ؕ�<�HyAG���+��������ҋ�A"�<��T��;o�~@C�ޔ§��LaQº�L�.�>f�c!'��n�k��0��q�T �C�o�&vp����Ղ�y��x�#���v�4��}�1�W5�!Bvm����֏k
�S[�3'$H��/n�5ꙝ�����/]�".�*���q��X� ]����#�7�~��a�k�g�e��2DI��C�-/c��($˓A[.2X�6�"��x��|%��J��sw��"'�=��O��D�4QE&�\�y4��qi����Oȹז��^���m�Qm��(�_���F�MX��.��d��a��=����Ե�o\��`���<��:��:���Ĝ�υ�����G&!���1ʸ8��/X�]�jl}^D�w촍׶�Vd�M��P&3"���kJ2g01&���c�G ��/�Sv�*�`�3��)����.�c|+I<LL꧟
��W�����Ʉ�%��]jȳ�*S�'!�s��+�볳KC�O�,q`H���P�l���^��9�˛��X��<���8Ի�čǞ����4�-)�[�m���i��A �����G�?}Nw;t��/͈�B�� #����F�l���d���cFd#i3��Z[��!���PW=&%D�{�|N:�[�˻^�i��ڈƠ��T.�nN�͇Ba��U&26aRN�\���� '�	��NG�[y�=O�fx�j0X�D���A��������x408���y".*m��$d���:Fz���iYF���>P&�g&�D������� ���͌(�s�1:�l�j^��$$OO�[�z�j�}���7�ٲ~܂�|�^��u�;*e���Z�*�h���+z�V���$ܠǡ'���5��Ў_iYLjE�ZS/XoL��+\�A�^��fA|Ia�H�,��?&�=D���O����ln�Ing�:ߋ�K�O��)�#�`�`p11�t��\�0=�ɚ��&�P(�E2���7c!��5�c(�"NԳ�|�:�����`Тd�0V�J���s=����$�8�.��F-�R�#��oT�E��X�X��ʟ���p��}F'�%Lw�UK�[�'�p� ���]i2o������]���@{׊����"��W��G<ۥh�=�NK�����WUX��5&����8�8~O	t&�lͰ66�J<������ĉ�pI}��So�K.H��d�l�=n�X����(s�׫N��GƮ��������-
�����_H��EY�z��}@��@��Bq�6Mv'��yorH�$?��	!�G}�e��` �A�P:I�<�t*{�W��)����
!�g�y��
�	Bq�w5p~'�������ژ�2�����w����Whe��4����a���W��A4�_}���);rE$T>P��:�j��W�>�|5�n�]�ʼ�'��%>}�"�	�u�$<MK�,Њb�rv���ŷ�����78\�1eo'����Z�"�����#P���Rtn�I!�]R����n��eK���Wo�n�EJL�P#�4	�bj�"�l9"?4#��o�����8.^��g�j[QLE�]vϪ&ȼo�c��$"��f�����;�{;�|*O䆮�b�Fr�Z_d��wpF��3���;&�O��/K�X�[��/�\f���>]Ɋs)��9�7*�����W�fSB�˰���?�<z,O��������[ID:��[�!�"&-�ié���yڷ��ü4:��Np?~9P�ʍ���ꅿ5�?��T��\v�u�}6�̇�&Ӛ��~��	3(������+یH0�g��eؽKd���ԭ��\�1`�0����I����Y%?�utƪ�UıJy��C�0�.��E/#�nE's���+�6ܚ/�H�bĚUN6A3�\a��{ba+?��3L�ފ��6X�*�9��p��11E����OCiD��u����Ck�y����o�)^��������xI��z+�2W� ���c��
���P��K�7	�
�����	gcɥBl��N^K3ҾǷ���A���O	�QQ0����zBV�=}��Ԩ�ǰ ��p��_�g*fR�N���?ǎٓ5�EJƚ�t���w�
�3�~}��&<�{t�s �i�򄕲N���D���ӌ�c ��/#}��|���"�99��o�GCz�g��[ su.���ao{y�ao?���F�F&�^N�������jE�� �7]�/���9eB8����N�D �S[�O�&d���S�}���cJPl-�����&\\7�e�H�!���{��I�_��(�A�ʒ���m�Eo�-NGg�����h��X)�e"��v�����m'�UT���F�k.�mI�:>#&Cm��F>�̥�n,܎�9�!t|��K�k6�T��,N���=���:d%ͩ5Fݮ� �g݃����AC��!L�Y��u�؊�T�+,R��'x���Ԍ�I���u؉��	�.��6�GN�W�T�=�^�F�t����ق�~�ן9\�����P�@gl��'��=t9��f�dp�]W�����G!XZ�n�g!�|�5��9�C�|�
��n�����Ԏ��!������Kg�����XqR�R������"��j�Y�QQ��	X{�\����x@+mY|��PR��X�]\�{����x��XO�(�䘗C�y��Ni����.�h�����c��gc�����ݕ��֩e�4���~�ei �=�IR0�F�Q��H�_4!��Y�4��� ��X�ޯ'"�bP�Ӷϲ1���%-��ѐ�*�|�"ꩦ���2�Td��>��J�����c����F�v��;h�)σF([G��L�uv��%Dm#skK�
�b�Z"T�HH����_3^���yH��\�����4B�[����ʸ��8@����5��Wv�����#)MZ��ݨv"m������I����AmG	%�������=�0R�g�d�� գ�j,��(D\4�f����â@���m��5�Sv���bIS�SE�w[���I��#��xy":Ѹ��^Н����	c7�4��;��h錳��&d�`��Ȣ�Rе#�IC[E���1��b;�Ѳƈ)5L�>s��os�w/7�ClN�&ط� �^`BK�q�w1�x��J�;�nX��r;�˗4�/��t'��D�tr*�|����3Yj[sa �s�ڼK��O���D�6ڜ���֥e<b��\êX�_�2�[U��ї|Pg]¡'�(Z(q�,v �O�"�Mb)�5��3'��AOb<���\L/eK�H� ȼR7{�ժ-;�(ې=�����zY�-�v��D	��IV.ebS���$��ѷ�"@"��W��[o�p�������pa$D�F�l������$v�.��~l�z
��P��ύx �ߔԩch�חׅ��B�J�}�v�:*'FU۽jR�/b��01,(,vÌ񷁛�I���-�3ˣ�h4�5f ����I�/]�zL�U�P[�i#Vf��_&�>�?�l�aͶJJ��T�%X?������A�G���0�2���`�����pT� �[r��k����� k���o��U�J���_u��7�.�2��F�!.�^����e���D�ZC������7�Z,�?J�u��8����A����ߣ �XfF`��}�#�ܤLDvf _[桗?��Lx+�B�x��A�>|�-垭�E���U{Y]�& B�?M������k�ň��Gx�cC�a�QYJ���%�uAU�;�E���IJ)�#�L�Eٸ��]Շ��� ��Y�Q78��\o����9ϭqsiH׫��%���4J�S�����{����fO�{6-�W���W�pũ���/�p`���0z��Kl����X)	:��`w�JѦ����������W�͠%Km"um�[v]>����?!�F�P8W����d���N�К�e����n@-Q#�C�LT�0���B+1.
�v6�!�;(�l$��Nx�R�L�wr�d� =Ʈ���Hh��F�4R-F	Q�!��&��[�s9bT2�wzCDgbb:	����<�̟ƿ��Z�ɢ{'�ː��KF[#��ORܬ�2�����m�Yy�	ۣ����������l(�k2L�,�i�^�:Z��	'{���#(�>�&���e�Eǩ�L��a��N���mt�����]��r����CU�	�P�hG��
��[e9_�C̭ÙM~�[��m�������vU�֝m�'�$V�?�KP�sh���P���������:��N�D���Z�K3���a�N]��r�!D�Q�x�їH߷��.|�-��V�{�"d���C��R�<�-`D�ܦ���_�5� �����eZ�����2N�{��2]��GW�ĄX^�<����4ˋː6��6~�o��m���*�G;�w���
�\:��^F���G1�
X���*�����
�tRK
J��#�v�s}����aͮ�����i��P�f��R�p������x��Wr�ļ_|�����¼y\] 	����N��Y������<?��'�e�-�ؑ���r=�����H�
4�e2M�c�_�܃��.�)R��wM�eCTfk�:���?v���&��ҦW%�+�� �V�M�������%iy)	�/���9Jއj��+@a ����f� ��%��a�S�S�0J�A4���b���&���?�=����
5qA�ڋ���ZN 4���S�j��;���������T���R'�
��q�x�g���"�/oԄ(*3�<(O���
`�)\ُ�z�)	��_�Xu�y�>G���ڜ�(D����h]j�P�x=�������=$qq��IX���Vt&*�oEQ�;���=���b`<�=��bh s�LJ��`�����-���z�<΢���
 e��l�ޮxd�TU�����1_�@���L��k7�n��r�
��S�#�*3e@!�b��|�>m�ڹf��yR�H�!�94��5��4Qx��OʤP����������B\����f8�h%�Z}�UE�\.�9���䬘흑���iF3H\����ZQ�����S�⁴9�-��w�t4ux�1s��3��⭨�/��O�.��"�:��$S�
����c�A��bK���C8	���w��|��V�#i�}3���5�5p}S��u�4�&gV�y�G�!�t��T�����$3q�e�|)��wP-=�)ŤJ��ۡ�b��\@��A�,w��x��2�|֬�K���%�Ӱ��^����#�E��a�IW<�&�J���$WE�o.5��#.��t�I�R�-[:O�a���Qf���<]��8!�lA�{أ��͋�0e���@*V�2[;`��M��l��+�gz��\M�/n�~����kw�% ^H���O��F�e]���r� �ު�y�դ|�����64�0i��`�Ǝ�Л��D��OW�@*��r�a����K$uȼ0�	UMY�~�����#돹������R���C4�ǫ�̃K]
� ��7�I>��a��u��n�,�������u�K�� j�/]�t�Y7 -�s��Ꭲn�����Da0�1 {�4+k���\B}�Me(��78�z�y�!����M��` ��д����)��레Q�4�k
���3�ܠB�W`u-�,h��̖Đ�kF�0���wn/�'�參$'���>2����4�������bZ�j����w.���d��jͭC<��<U���}��@tN��x}��<џ�a,�M��V�LV|[��~+R=��,}��ʔ��ь����_�)V��ߣ^�-N^a�c��a����Ӣ&�B�$L����)-'H�V���%�Z�:��Q�۰�{���C���Ys��#��'�y}�
��Y��N�hLaGI�0ti`dd���&�faA�m�{>B�jɚ��[떭ـZ���|/d��!��5&���H�L� ,�3�������g�����yN�Ԭ|������u��.���k'.�J6O���U���A;`�Y��R���N2x�-�I���Ac#̨�ǭ�OH�7���oѽA)S�#���*ҩ�R��UB��l�4U	9�zݑ��Ug��v��k�`�y�D�ڀ����S�?���jD���jx���?.�
E~�\�X��w���<|vק�8Lq8q�߇��d���CWA�geRr��,z����wkۖWX����	{y�KZ�֙�~MA]Ө�����jxf
��S�TMU��z�[u�Ʈ��C_���]�#�寭z
/�/O?�a��x�����'rΡ^���E�`�خ��&\k�W|�ߩ8���< Ge�N�Cĳ!���U��� @�<{UX�?�W�h(v�;
��~b5x��8��\�,"�m�M���U��~l1)^�J�yBA��sM�����V���RE���[���^�dFt%���S�t��k~��>��E���{���{ /�jV�ϥ�yR
�P:��Q:B�~� ��+�1<OV6U@<��Ϙ�`c	z�('$H<u/j�Pnq5�)dX��^�V2)$K���2B��JI��S���
���+9�>P���)��'��V�z��l��e牯�:��1M�������h�qRd�Yh�*&"��*��Ӭo"]%�:�\��D�Myl�ٗ��6��;d �� �T	�ϲ���5��[0���8��ڕi�������uN�n��8I�8y��!= �%b��4�۔���U��d��t�6�UՓ�G@�'��%X�Ƙ_�t>w��;��d��=�!8�eA�8�Hh������]Y5b�pGGC�mj4�?�axda��~�A��{��WV�/	��Г��'�OU���_�*�E�k�T�#��^��gYb�g�T���ӭ�_v�����Qo��l�5��O�M���R�8�b�D�fgN��iQv�Xb���HҘy:_�����rU��ݳ�R��8�~�.��(�8���g�� �w��(e�2�JL�z:E�WO����zA���"<J����m��ß�Ho�����~��ap>�����3SF�z�1�.��9�
x�2�ܻfkd���F����H
�����p�O�2�I���	��v:�{RU��/�z�g����)��Ҁz~ks��2��8V�wu��h�HPU���6�n/��<�zV�vK��Hw���D�X�M�;Ul��=�?��^�~6<&�|:�k�h㙿�hs�'��_C�'?DT�����H~?"�v ���*nMU-@���Vr��ש��f�{����:�U��}"/�OѾ4�����*�#�x��VK�fԕ�����xC�7�6��͟ �ᡐTx�7��Ef�va?�y�-�9� ʅ��G����1��7Ĉ�\�U\�ON�ɖ�$+a�S��	Լ\��R��9��|��f5�K]�h�$�X���&�P6�%/��!��#���a4�,=�0��3I�88T"MkT0I�[������yݜ7
���U�z��_�6B6l2�w/��͓n��L��f?/�����U���L���X��E�P2y��?K��&)I[���T�_�gi�������0�҈���t�kH����FCл�<�¥������z{�ʉX*�?U��)
�ARt-�m�� �U�d���*�tTw� ��tZ�6����1���a�v �L�F"(�-�u��ޏBF� ��5ģ�A��������|��`6�d���mt}p��5�,sq������@M��v�s�|��P��L�c��B®�S ��X��h6�:�A�cR��:@m wF�)�����#�L�	���Jyמww�PB���Noi�}�q;�e�ws�rNC��}Ud�Mɔ9t:�Kt	��滔XY�"O�S	��D(�T��B�m�j��U���v����7��Û��D�yÆrE	����ukT�����?
�^M�b�U<ФP�S�͍?x�&l��Cߏ��_��}�/CtO7SF��}�Uڵ/e����8���"Elͺ9�~+U�C��D5��Z������]���)H�da�� [��S��+�	ϋ6�D^bz0��[�"-f�8����"�V�L��\��f����5'J4�8_	6�&-�:L���<!��,&��]i:���ӓ>�nڴI��m����+7��� ���Jv�6S_�B�D�2Iog�	�13�б*ӫe�������t��2�c�}��Cx�!/ϳ���>]���t^�3 �S�(�q�[z����ʥq���c��arGtq��`$F����v5jJ�KȎ\*���r���e���W-z�ݩ�#�^`8�yڰ���x/�cg(�nY%潅���� ���� ��&Ϲjw�	��{_�O�ǁ��<�r���4d�ra��I��K��DS=�8R�I�ވ� �y��c�i���� �E�1�(�����'H�I�#�̩'�k��x������.�̂ �ɶ�SYL��no-^\��|hS_�N�G䯐K��b�%�lUxS�3����L��؀�GثZlc�-��1̼B�4@j!Ps"X	�	��!Fqp���_�6�&)��y�\M2S��a���b��<3�d���yF���ER)���@Y�`IbP�AY`_��Q��M+��Alֺ/k���4��  w��������F�N�m{zd��O�����^��nl��	ňʶ%��[7����_� *���]p�E�nl�2"&�����ۥ�$L�(�w�y�����F�%ӑ�ed�u;�4/VSm�Ǣ2k�>�g)���7��!������8Q�W��g�6��M��(��$��4�o��߀8�3�uR�c�C��XA	=拮�  �4	���1���l����OȨZp[���l�^��3-���b7߄�*k���۪�ܔ���t��y����臩�}��o �k� X	���(�?��$4�gM�z\����I1���C����MQ��pN�j�ڷ�-���ON����/�['P���1�3jX��i6/�Pt\����%�\h����br0S��
�-��?�j~�����,ͤ?2uY<���.� �_��+>�2�Қ3.{B�̓W�����)�V8�>b_���MGP7)��w�u_CV񣵭��}���d�Y����M���Ɛ���31;{}W��Z�;�z�Q���A� �	.A��C��l�wz�tw{?1o^Ƅ �b��m�yyK�J�N�>�g�
�`��"�P>wD�WX/���yv5�e���4b_�z8*�Gӑ�3v1��Tw!����t�k�s�L�y�cI�;f�20 ��`d�v�
�l�初���hX~S�b�O�m"�~�����Xǀ]��H��1�s��S:��:^�_�U��Ӻ���gيv�09[���m���?�pCD�X�X�οԄ�x8�~� �~�(Y��l�p�J���zB?.
�W}I����W.~n7��p�0�RF��w�e���
�q�}&t�ko�7����H�=&������!x�kc7�9�#��A�jӀ9�[U�^�ly�-J��"�c^�5w�1�J'S��&Mkߗ�s$c��	��A՟��CѦ���͙��BmtrK�uF����*�?iCA�/���8�Yپ0) �x^��07G�U�V����]�~?V47��Ō��!f�M��ҽ�`:����,q?uh�0_��3�fY�tI3�O�S�D�K�5�_�:|ݟ@h�?R=��^��]´+t4r.M*�DZ�r_�b_kz`���t�"��GxU�)y�
ub.+Qsb�_g�
f�y��LZ���h�;��Y�}�Q��ƣ�Q�W)��Y9&|͢�w��Ød9�K�zW�"�T�f���(]�1�*����4E���Hw�k(0�`?*���j�83�S�f# e�<N��v3U&Qj�|yɿ�U��Qwd?������wT��6Ajy�]�>'��
��e$���e��"Ie�k��|��%��jZ�yA�8��!���}��u��mS��Jm�q��=B��#��T��c��#����r?��K�0@�:zy�R,t^��kU�U���d	ѳ�Q�&��*1=�H7A�:�Nb�d>��-O�9"��vBA�h}�*�l�A6�!�V��ޣ�^C��G�u2ER2��dd2d�$g�CԿTqƜ=�~=�Fzє�x�+�}�+*���H6�ȴ��n�	~d6���mV����7U�	��th���$0L ��N�q�_/�r,h�&�c:
_�"��{�ǻ���Rd��-A���`������� �-\�V��[�\�0,��.�q(��1���� d��%��>��*��b�g��z�R�J�Y�S�i�E�~0��S�*�����V~�_f�Uy�f��/!�����K�x��h��Gf8�K��fM.˼�`uq���E�m���|�=?[�{ag��KpU~�Y��=6�����W(	������hhg�&E���*9�ʆ�%�(�������W>�����Od�
���p�x�����'0B>0���z�0�"�)Jی��v��k���:�`�`Z�����k��
5��'l��^H�ƞ!����
e�9߻Z�9���5D^�k�MQM�hW)�r�ޝ�!:n^�Ɲ��@D�"�ZV���"�̏#���AT4��͆+]��� �Jvˈ���i׺e�ߎ��otn�C]�'�$'_e~V\aS�V����Wv�j��@�E��s1�O]���q�t���ٷ�(��
�� ��b�����D��Fv|�̫w�,:���ǉ�xj&0���"���$���QE9����ɧtk�u!�t%�mh���mP�͹F��c_{p�$ߐ\8�۾�G�a�@$��'��%r;�G�vɷ�4�|k@�{�֟t�Wi�JQ5��<���J%<*Yr	�y����;\�&A���N��v��U��.���/&�^���#�JQ.��ԝ���
<�w���d���/y/���#����k:%���g���e��V���{#�9��F�17�$�Y �^\�n������CQ���Ed���J��c�q�1�z('Cmj{_��x��'Uu@�E��d�|@XL�/���I�ޓd8��V^l�	Y�D�V�-F'uxw�nl��-�yi��,ѐ	���@7�@^��+�� ɞL��
���-���F�yF�v/rص�{#�'SR�حM�'����0�°Bˮ���g^����0������]K+j�~�����q0�dlP��%2eM�"�P�C/�@���%� l��at9��ӳ���· \�}Ŷz�}4�$:�������!4�]�C_�#DX�u7�U�6&�B�8�������
��eg1V�5j�w�_�К	a���$	?�����S���,�R��[�ӞyO�?ϱ��(�f��z�,K�%���4�R�f}�d閂�p;fx�w��46��O��;_�*����$HlI�����;�IZ���V�h?����,�Vv�!sk`�����l�˰Ai�z���k'��"�õ_`G�;~�mYO��e��(���%6n�z���?gۃV�2ތ{�Gq��H�ˀ��TtϽ�e.�-��8��d8(�� �~C��$�X��� ���$��}�����n���	
�C�� �D� ����Z�����;i���!LW���2��剎R�D��b5��ܱ�3�{8��Kx�)��]a��s��y�[����T{jac搾��b�I�q��[qxV�wNIT� �?;�ɻ�-8ȓ��
8��[���@�g��z~W�}���`�����`����Kyv�[����' � ��f���c�#U:f�C�7/ԜY���+�HQ��g�q��ح��x��=�}$z�P���Ǯ~k�r8��z{�U�\F$+�8�������)���"�Ѭ�r�� $���}�F^-F��x9�;6�1 <X����OxEWzS$+>fTNbW0^�8,@�;p���i�c~�h('�Li]eȢ����4������]��m9cC�F/��V����v�(С ���	l�s�44H�!QڧP�~KI�E�v��o��!����=s� �>���<���?!��buZkFX�cJ�g_'����cd+]_��LnY�ezT���l�B�i��������#e��9U'}K4��M��zM�K��@�V��E�G�
�1 f�F���C����݉��8�G�%$N�G����R��w؝�4j�I�w�5봷7Q�-���B���'ڐ�G�w�R�E�-X�����?4���G m������DH��0�C�����ٝ�Cmpv�Qf�BQ���F����Ngu�u-�>�t�̃�{/�Ҋ�L��$d��Xg'�cP�{�������aܹ*`8T�VO#�m��+����<ۦ$ߢ�����=�GY$�veǌ@ܹ�ڙL~T0�Q��I��X�%i��Zm�����?X�VTe�3X_�~ב��RP��1t���p�����y�.�����a&��|]�)qK�?����z`P!������`	�퟽�Ƥ����x�0���Fd�V�R�]ޓ�]P:���vz
��֕�s\�BC�ɼ�����4,׭�Ϟ�����ƈJ��p��3�Ƽ������ 6!ll��&��.�|TB*8ny�P�~t���@�<��_����Ь{ծ����JP<�B)h�-7���"��p������&a8�s��񁱾B�Ȃ򃳌?��k�c�����AK�[��~B�Ǔ�%s�v���+��s00d��U��/��qq@₝r-��gF
,��"�a�V�7�8�T Wo��ʵ�PK�I"�|�r@8��$:5����]*���X��"�����<��j�vd�--�����3ͨ�DY�����}RK �v��gwL���;��R�jjfj
\����[��(oK���h�koĀ�$`,�F��B��N?���'%�Q��΢�}�!��f+�����X@/�@���΍�N�3۽�9[v�'�t㓱SUIU~{�)L�ɔna�ɮ�=~�9�՗��+��r'^Am�P��-���U$�O1����B����t�ҏTw��B"��������wf�,���\nɢs<�LyDu�@'�Fa���ow�/νW�\��NSZ���\�em�X�~�,�����6�ZK��H�MXD̦�>�
�[���9e�َf���>\��ޠ'�b9.j&_�d���V�k�ߑaDG�"XLh)O@����)}�K`~�:��Pgo�=� �/�T�IWc|�� Q�ek>\���(߁!.�5�q��6���#
T��JU�Mu&ac+��l��US��=WC��������O�hS��kCX:[z'U��T~$���p܍��%0+�OTF���*�f�����0�?��Ζ�����鯨BV��R� �����u
	�o�A0`3Lb�\OTc���z&�MqP�ȩd�R�ʿ�_aN�%�*�s�&P?'��/27?��׮ũd�Q�l�滋7�h"/�"Mw��HsJʥ��y��%�� .4 zD �m�:�4(���w
aw����a���!?7Ƞ�y]��03%�>�;*�D��f�wW�fp��N�5�ޒ���*��k�8?�w�����
M��Q$�7�����Ʀ��m�55��AOX���XyŠ,��"����8+-�O�?#`5����g��1�Vl���{+~*�����*� w��-m�3�Ǧ۽�t�#���c҇���q-�n��v��J��̦�%�'���g�[3���USZ���R�Yh&1� �B�xm��~i��:�ISNXra�}4�/]��Qjr�5�E�ȿQ=�'ꎙ(�e�,� �K۞�Kl����T1Ƿ$3�IH|E_�@w�ۇe�g���$9Oխ�^OU3�׾����6U�jqj΋R�㛞d(#����Jl�kڮ�ڃˋbA����֥������ĞE��J��4&�A�8�VM�C�����|��SV�P�����=/���@��)Y���0��%g�1�Ϯ{�6}N7(��"�V�]q�'�W�8�ǊVF�	t�@�n;���An4���q�Ii6 ?~�2Ľ$orLo�6WA����07��b��@/s������|�in�\�~�m�,��͛h��]��rZ�F�b	���w*q������Lu��W�	6����CM�Iet93�v����@����X��4�{�ngN�![��	%3�ܖ���W�T����ZY�|�K&I_�G9�U�%P;��)6?.^��WWȤ��#��^��d�aˤ!��)��_���J=6TG�ӱ$2H���;��t��s]o8�2�I��aM�R�n����e��� py2�bq����5�?T�EH��t�]c3�h͎v�:n�
`��)�n��a�+�|��g��iR�򹡹(�s��?�Bm�},A��:�[�I���GOE��X*׮	����䪇Tք`D(ܽ�`al+�7�����`%hpU�x~��8���lmL0f��e<+_�W���W&8���������h�'>��P-^p0)��Y�u�3+o
ym ��}׀�����v��m]7FlFH�w��@���!L�O��x��,��%�߽U������ �����c�U�l3������"˖�"�IG�=lH!-����#c(���yȼP;HَC�f�ƍ��/X�Ģޤ��1�[I,ľ%���Y��kN�݂[�#}�0P���7��%���8�#����OT;ܓR81}5��>TE�m �1�pZou��Z���uKv���,�3�$�%j���]��.�@G#�Xx���?�c� Ӿ�![�c���c�ze2�Y�+P��\�,мm��b�a=�V�JF�����U8��y*hY��I$fƉ~q��\�v�Buk�����I����
�`�������+�'ъ�{������ו%4���KD�|�P�~xs0��%���\��e��f?*^=��$���w>{?{M�<أy��9w�|fH<6Q?��e����+.YL�X�n8<k�,z=_�p>�d��/����g)���|����F��I�%9��,)>��3���p&Zza��`�&�q�,T�ApX�Q�%��9c?���� v1Q���dk���M΀� o�!0]�H�-�ӺK4�0���F㘶dK�@E?�4��,C��I�|;�D�ϩV +��ahG6.NTVy6=ҽ���Y.�xT�#8<��X$�U�xB�{9�t�����s.2h|Z4�|$�q��y���	�p��\2�ϳ"hE��PjB�V��<�Aߝ)js�:l#�5��,���)����;�v�݅���3��0�Z<�b���d��ǐQg��~�\�C�&�~x��]����H�yp�\�p.���:S��������H����壋hKa��8�	���5��%�VU��y�J<s���3X�RS����%�#Vz�I��;$24+_c���҄wވ����(���L�(��b�vŶ*iT|fـ�8�Y���(s�M5��V��W��֏2=���iF���ǃ�S��=���Jq��ټ����A�������9��솖��[%O�(i� #ڹ�=Yɡ�r�s�qg���k3(��e���˿	���g^YK� Fɇ�(j�qb���'IY����eI�u�zt���"m�I<�3d���Ƃdh����]?f�A�$�TVtf�5��pڟ�x���4��7t5���d٤���5�a���N�G�WN�$�%K��aާ�$R�I��o��1
��{}^�{�����*�p"M��:����b<V%���e7���p}s;~c��ۉ�+mu�a@�U����\��?w�$����/�v����Nj�F�9�kQ�l��L"�������W�1Uu��̳�o�mg�B��;�_�E�d�����ϵt�is���1oɀ!�b���b.rͰ����⾤⅙�sl�Zx�����0��,}zںЍ�N�\��{��6�5 ?�P�]p���׳4[�T���t���Ĺ���mH�� +4�� ����vl��/	S����~�}��[��ur Z.�g��\�;2w�{'ki��ܝ�
k��V�k�t�wu��VZ�_����PN��.Ѳy=g�RV�)J����<@R�z�������]��,ԪݚN^�x��V��}����*�.+����
m���Ոt�'vz[sD���`�	D��{���|���D|�2�c`;���$b��!��E�V���������#!��M��mq�uG����ܪ�ł��? �T9I?ݔ�X]�\���x���j��BI��V�3&�Z;O�`�:��t��G�����xp�Қʶݒ��?�ϛ���狩���T ���E���_���?ݛ�<�OV�%��
z�u�;�	C��$���ʨi�A�8�ጟ��0[q�ZM��j1�rٻ�m0�dF<	j-�HZ>H�ϓ�������UO�p��ſ�W�,��q	�Ƕ�6z�ͻk��l-'��>3R*2Z���{�W/|���9��A!�;��j;��Q�Ñ�4V��W���{E�b�C�4eL`�٭�+�ph��(Nڗ�C�����h�S� ��
f��a�ޚP��ŇE.#�?�3���������+-iW�ӧ��\_F%5�:{܌iQʺ�~�l
ȴ�m�	k�#�����6��zS4�kZ�Q0abОr�:�8��|!��M�N��0�x�h�|��-�ވrL��c+�Ѫ�;q4�������N�Y3�M����A�-�c�&])���h~6�ܿ��ȅ��(\M�t��
a�5$]:v�i* �:/cf B%���*m6��U��c�8I�0H����7ey�
l�4"0�!�]�_ɔ3�(z8����%������*�o�.��V�sT�������`�OW� �"'�R;.�C.����K0r�V�rU<\,r��Ė�|�$�З3���#�'؟�"�VPV9%9�@P�z�(��3���/8� ��숃)�i�/5��Q@��RU��v�&���D"���%<�ڵش�{hbxğ%#>M%���ܵ�&���4؏YB���1��Dy9nJt㦱K�\��n���Q�5�G-��lj[&��ow�G�"��M�F�|�O/h)��pλ�:ߨ�9��\b� 9}�h���5�p�����/�4S ��`xF�y�;�Rn$bE��J�䃮��C��H�� ��x8�u����vB���q�%�X9���F��PJ��ܩ6L߳s�Ϝͅ����p�v�(.
o�4�N��屈���.l�Z7��zݖ�w(��qA6)����nb��SM�RlO�.������P�ϲq6�Cs�|�m�0��~1A�7-Wk��
-Aa(�$�tN�rd�}ΰ��&UB�*��+�e��RaOp��+u���:�>�<�*;)���F�+=:{@�:�a��(�h ���&)�;�����@�yw�K�Ё��V�����=btT/�2�D�8u��4]���6r�}�N<�������#����rF9	',�oαד#$Օ�X���ը��Xb����M������;W51Y6��p��9�$*b���{�i��h/�:JY�Azކp|כ���^�_�Z��\�^oY����R���*�^��)���E�� �	!�?�;""�@���X��@Ml���nv��!�m_E���w�D�u>�5���65S����/|b�E��V%T�L��*�$�.��6�%�ywD+{��4�$�G���&��6����:=]"5��|G�砳�k\���?:t�r�zY����F��J��X[R�i?r�TƵ�:��3%d�� �n��jk�*��ѽ�W��\t�t�����UZ۳D��p iog+���/� c;�cܼ�0�N4���~���y���w������)�_�b�`e�i�Q���+!4�G!|�+<�Qhj��,s>���,-BY�m/a3���6&	n;��0N;nN�R�8��@K#��l�������X���֭�;otx�N(���D�9y$Q��� ��V�Hc�j�<&��y�_rkM�	����+>��	M��op�:+ 0��UQhui�׶-�Z���Y$�2�g<j�<��6�fp
��+e��ۗ�Z�9��ܺ����mڣ��Xߨ �
�w�x���Qu�>�V.�"�.Ɏb^�9d�Diu�,B_���Bw� �~	 �>�F��ePU�I0��.��L�r�i�7���I�A�M�)��C
[~�Qt�=���&K� 8}���'\"�->P1�Vgn@[���r��|;Z�9�	- �hV=߁����*ʒ�U���)��ׇ�´���Q���>�����dQ��d�D&�uw��8��)�p��ڝ�#��!���P�j�v�"�c/Z����W���C�_�t[��}%�
����,���90�3���M z�W�/<HL�B�O�������o�������YOA*pn"��YZU+_L�M�5�~���T�o7�F���`���!�rz4y���o��aV\�wk��/�-5�ɦ3����R1>���L�.��4���'��5{,N�3�LS�Ȃuԡ.��~�*�qj�@h�CyC�D��8mT���[ᝡZ<DE�=�
���+zQ��8@�B71�&6��Z�c;IJ
:��K�#���{��2#�{����{Q�f�������
L�Cl���(�@����8�/?y3q;7�#u�� ��ȕ��E�����47�O*���S�A��n�|.	X�˞�҄j$�F>�Z��#`��Ǣm����վ"{�6w�S���a7�}M>i��J(�RY��(U �� _��P��PE���#�(�h����<~F�ۛ�0���0��6�-�HV�G%bf$u)��;ʌ�=�#xx�W��6w!�0	���?U�JM�F���J�Oq�f�	����5����?4#���ɝ'��pn<�>�s˟op�W��>�ў܂��e���1��j@�E?*�d�@��z��Xϑ�]%^ �t��o+������5�+eHq��ɽ�[TߠKN=�A�2���RIr�J�F|��]�U�	^0�,l+�ɱD��ύ�jm���ϡ.�6�8>��ǿ޽p_��@&��{?2ѩ�Gx�2c�c�q��E*7m�d�幌�+|��&�����K*���)�@��W��?�s�� $������xAXE\R+%p�>��R�Սw'~���$����5pW҂<!�S��(r������d�9<�}�K���!��*䒜A�]�z#�'"V.I�P��yMϏE6YS�m;?M����=���������Y�sKv¦���mGY�o8f��dnί���f�W;п�SEE��4}{.�!���;�a[���ۥ�0ӯ�<d(|�Q��#�#,�ػ�_�>j���؃�V���N�t#kR�U��.'�7��e$rR���B��NE��S:�N{3m�&�Q�@:��>=W2*��}\�mNmi�j�a��}~J��y3 ���/p�M���/$�}���(O{���M੷����٪tS�T�͜�s�����&%7ʶf
-�>�Iƴ`A��k/��@��s]')��~{�a�����)UE��+���q
zpu[��"	�nZ�)����U�3tE~�K"7��k!N,B�..>���Lvn�|�ǹUPl�0����A�i%�K���)�������p� x�I���zh�
"JyT��^<�����sY�q.��D�a� $�nt��qa8���V��a��6��$'��u//ډ��4`����-N����X^6�b��n�C
�&:�~�܋yB��} Cל��pĶ. B鹱X�S�Ƶ��z��1߫?��nA�q/1�����fp�V�e�s�q��KR����ݹ:�>3H^�<�fUӨ�lcm��R��&P��LN=]�S��4!��k���P��qN����d�Bv�E�f�꽃Z������1��T��J��3�-F�.wm�/�A^��X�J�^�v=�z����V^q;��.���'*R����5ct�����ي���b�ȣ��=>����++�,��D3�M��~8%���\9��	1@-��U�e�4S_䱆H���:�o�u��:�W�b�'�}[CƻJ
�̀�B�",O1'��K4�-�9���R�����T�#���8)�hF��*K01�0�?9�N�,^��a�[P0Ή�~�l��
�mXtfX��:o-٪�#��&��/�Gb�IP��zn;����X��e;�S��
| �R�L_B����Lؤx�RZ͉�+�v�� ��K��(�\Կ�`������y�=�Z靧$��h^$���bѺo�e��0pO0{�	�o3�j���\�Da}�ռΡېg��K@p�F�z����ʃC8�d��kk�х#�`!���` �4	����Mͻ�a��AyǱ���bm��/O�G�Z�~���?ysc�n4�U�&�JMf�^= 7�}������=�ҹ���o
(��_ ��ii�O�`����Z�7�#B�?��V�y�7��t�p�yM���Ϭ���\fz�� jp�\���n�Bqh�㕽��ͧn��zT�ϔ����2�PV��za\����0���@����ò��"�[&��Y�&z"wd�a�Lܢo���X�=q�y5H��@�[���e�!Q�W�)���.�U�2���Ҹ�����Hu[�(G�@3ڤ����وx��Z�-�ٚ��#_q�u܂���{�Д@��MU �ALd.�6%<�_�,Ì�ָ0�p���5������4g�<�J[�� z�[v
$�?�a� �ȂCrJcj�3��=�@�o�#�)���Ro㖍�m���Ne�����5�R#eZ-[��{��
��a��2~��f�)�lt���-}Zc�M�������m��Ϯ(CB-�XC�{��Ա��ԭ�ͫF�����Ӗ�\�	����X",&�_��:l݆3v�7;.�$Ł@q=1���� �ϫ��%2oJv�I��l��9z�j�<`�:8�>�?KomRFD*x>�a���^���C8C���z�%}��x���#��~�_<��g!�I{,լV�)�|UǱ�T��`��_E�_�Irţ���k����o�9*�l&�]h
CΦ�t~W�3V�t�`��q�1���f����|0s+IB2v�	Z��2�,��Ĩj����	���'�" mܼ$hx����A��j0��qQ/&M6�r���h44f!�R�tFn���7�yQ�*J��.��Ͻ�/ܟ]h��b�;l������AAO�!�Kd55G�c抱D��vXw�k�3"�S�̀�M��*�g�븒$��gT��mU���aSR��z��Eyn�_���A��F��R�z��2��Y6�\(�Y�:�)w9�H�WJ���ǐU`Z3m��;ɥ�D�a�:��W.DHZ,8t6��P�i ����dߕ�m�!�q?)�D77�q�r���Y��R��6�]�Q0uݝ���-�����?�ix5n��6N��Ѩ��c�~��p�i����Fc�Ń��)���Y���1n,�%������J�-��`9�� Pjm����BQ���c�$�/,��bu�GR���B�>��f�5l�+h}:/��[C��)�y�c�brdHf�gYE]�c@�w���zB>�n}��/A�k�i3�e0�54�C�c�uh�>>���C��pV���j<��{hf[PF�@��z���L^�F����c��1��7���װ�
�j3FM��%�N_��H��;�T1y5�!e�e��n�|WHA1�$��&.[��ψ�g�/�A({#��XꂆXY��W�g"����ـSS��釃�l��
��g��:'�Ţ#��+��;����P�,>��8�D�3�W=m���e�j���%�Q���G�ğɦEl�C��[��@�g����q�-��f��J<�HE����sUm�]�2�����acC���SK[�g)��uD���3����l�ԡ{$^����V�e�z�:�pԎP�sC��Ľ��
�@��*��������珢lߗ�S�!q�b�]���1Ѽf���7F/%�`p��SR��3������\R�`�08��t��K�o%a����|g޾G���}��v��+P�5i�\B
Y��tOi��~v�&�tU'R��J�Pq�!���Q��(Ns^)>SC�%!�V������V�,�Q�������>ƚ��P��y��g*�+u�Pe[p��ރ�2��}IJ����|H����j��)q�/�R	!�B�oJ�|��E^C}c�V�k_~�ʋHs�j����I��G.�&'�y=}õQ$�(qA>�c�3S/8�������P���p���jӉu+������*}�	H���x� I������ rkTi�@�T��CË^4�Ӓ-(���@:�H �O��%�NtF�}��ە��=>���qv�C���S�����4G�0��B��FrjNnu���k�T?��H�11�䔤��PX��.N��ǗH�B-�-�J�P�J�(���pt�v�垻۠T���mɢ���QY�HO��KTO�ʵ]��a���P��W�z��$���YJ��]�7ǅ�8%�� �N�F�R�A�C�ϩpϯ�V�������[U|_HW��'�������P�f4��\c�J~h�6%4l�L��G?>���2�%C	0����6_-�{ڤ\x��a�	�i��� 1�ݰ�&Q/�����:1����m[�>J��02s�uδ0Kb��G��m��"S0�6��¹o��/�[ef�o��+�W�wv���n�J�
�M�<�ZW�3��astӳ��z8Ɵ��hآ�c�S�t�|�6�r����^J��:ٷ��Wn���Xx@���
��{�"� �ضJy�x�d�h�׆E&,O2��!!����<�B��G��Z����"�4g��tD1����� �����$�O��sO�,��`�!��Q�Q�����4L&�`8�}#�v��O����8/�d��c�P"��A�3�3t&k�@�1տ�=˜(}�/����s�z]��s���Mlo�
	�	�Q�KL{���X�'�9����x��S�H�L��3zU[�ӳ����5q��lђYi(�;��r�1�6���6�9bf�S���]��$�(��H�y��x�HY;R+21X�I�Z��R^��' �˚��x4l����W�q��V�+��:'{��,r�+�=�������O�3��)t�<��0�u��@<I�~.��seZ��%ο�qO�tl��1��C �f��b�b���~01�=�7K)x[;S�B�lc�A7&����IZ��T��7V"�亄�$��.�[J]�S��f�e�:�]T�h�W+� *'P;���5�a�5,gYZ�ά�K[JzB[��-��｜j�'� �Ý�d�k���f+�/����[B`�m~����-"r��̽p:W�J;y��ZB@QC�5p>��jm�bg���Gdޓ��Uj����d�� �k3�,�FQ{5G��0�������螑�b�p�6��!J^F �YIe��38�ݑも)'FEؘ�%~l4Nd�\F^D�d_����o���i{�5У��¦����Ǩ���b�l�zI���F�D�b�����B�)�#X-Wo�P�-�Sd���2��x��Y��ܫES�Nh�X��j!ֲɫ�%�Z�w��VxWf��Ta�Tfu��S�|�ÚG��w~y,>�����ī��6�C 8�����K�BUI1��p:���u��*�.�t��7����=�;�2zI���.*��Nw���B��N� ��]���P�G��RB�V�MX�2�*�I� 9�qR�
�l�Ud����:�=õd�	����q���+%�T+S�p`�bL:0�*��ؼ3a�d�L�A�ϫ�Lp�o9��KF��
�@+�^t�Z�J��׼���X��W��yс2�y�xF�0�+&IŘ<�d���o�Xl���Ј��^&ۖ�Y�I�E=n3���y���Y?��[ ������h�,��9�9��R�u�R�AA���~�i/A͙n}�3�ր�=_]����L���T�shk�)����aP@��\H�t6@}����D�8ʳ0̹q�4�������O5nw���ft�quNq�٦����"��Ɩx���A�q5��рπg��?��I��cj:N���C�F�)\:�a�����{�"�=^"p��q���'�1H��f��L�J㭊�E̶U���,�~�]�K�v��c��4��R�<c�}��0�r�
M�Ј��ʫВ|��yrJq�X���xsw u�+�Jf�9%�I�<�i��9`��q;-lv�����'�^�����ɓ��_��lߤVFXeg�BcP�Ҭ��xz�U5h+W�$��\!.�%3��ɳ@Uw��V����a$*��[�Qc�G��<�\���0��:�������!4Ş|����W������ԍjKۮ�wj� �]��,�ٱ�@�}=���~�ǅkUޥ�c�Q�����=���d1qb0�~~Q�vk�K�����L䗙�f�b'�p��bk$����;R%���N��b�@wfX�Td"ed�#��\v�m򬓔���q�<��nW�H������� ��T?���K�_�����3y&�OyΞщ�]��mR��(��.,��Aj�Yߗ�
��<֤�]��v?_��_�Cx n��p�E��g&�-�1��X�~�	sB��<���=ľ��"�"N��ڂ�v�L��f�ǲ3����i�E���'P�X�P&��f&�\�}yj����?��ag굠�3tón��<A8@R�ZS[ҧ-��|���f���}Ac��������;�_�Nf?�3�p��cd��K���A�rO87��:Y��<Kӧn�$���
�>c^[�Ѿ��Im�����b�j�~5�慝�˙���u��7�~A�H��\I���w�v$�{��=T�E���1
�TG!�)= |�t+�����/�J2ίK"w��7a l�q��b��(�6���֚��&3D �I�h�b�����0�����T��6ɭ����������C��w���~X��Mq]��X��Wv�Z���:�ѕ\����;�91�n�*P�;�۬�!�~t�C�� �jʥ$�Jt·i�Y��x�s?i�c!�x�a�?R��R�!�]7�5�}����ƒ��`�h�?c)�9UŨ������Z̰�]z�a��������D�G�_D���{��m�x�L�`M�Pl�ho&ؘ�5��HVEvݺ�`���L������&A�~��$�̔џ��0w�FPQ��&�`k�ix��D�?�s��I�Vܑ�ig����� ��D�����Ô,�l�mytg�U�ZB�S��ݴ�݃o6s,mV��;�Kw9��
����J��`���"o�K���@ȭ,���uR���?�mINr��<a�l�7��0Q�����
������󻞟��Uݺ!c�9�L4�C��8�ϵ�$'hp�B�Y���.t��\zu`0*��kק���V���b
.�?�_a��3Á��78�A���`b"O���
@��q$���/6��M[g�� �c�fZ!��ǵ��J!o��B��G�"~/���
�a�H��;�F��H��]m�q���R8W(�M����)�+�%�Y�z�c��J�!�q������E���>œ=F�C5�6�Gd��N�����HJ��T*x54�ɠ�q�ȁ�N=�����J�G��^��kI_��w���.F��i<�ġ�)f�p|:���0X�Mm����X�c��W�3�z'#�P�/��]]�Cx.�.4,cE����!�s����+�=�1P&(1R�֢��Z,��U��)�v,�R��"?�Z�Ey䛠�yZ�[�i4M�w���d(�|Pj@:�´B����KU�k���"u�FNe�e�?�'� �g���̞�[m�j�Y����?=�<�X���&��H�d��ҕ��X
��	)V��ǅn��x"#c��h���$I�;�J���olJ��5���>�JF���w�J���Ʌܿ�6?����2�qڟ�k5�'S���<Mhf����`:�룅$�z�#(I��=�XN�?'��{V^^{|y����6#�%�^KG�'�{
�Fo�ӷ�ݙ�NF5���CHh��4\x ����j35u�����c����t�=�5y=�GgCe���c���=m'�77��˦��F(�Bf姅Kp[{:�E���e%��O���{�������'AtP:ް<&��̅C�r$��0��n�6ޔ�-�}���숌͟M��)-,���^T��u�oap�S}oD���jp�����Y��[��	�ޒ��z+�Y- ]�k��fs�B�����BZ����M�XQ���D3J��s������n�w`\��*�j��9���1�]��%����=2��\�����)%��4o^U*���6�%v�$r�Y33ޏ1(���N������W�V�����1���NX�y/d��āU�p]+�Omw�f��Ou�f	����D>�������Z�eVl6х�,w������A�\	���:�X�ED�:}�O;�M�B|�V��Њ�����D���yD��Y��k��##�����-�oEQ{
T����|���ׇ�\�������a��Y�O�9J��Q��"%�vy(����Y=�C<��@"w�xbB���X4	�i�ap(�OZ�j2���J�TG愄r|���N��n4�ha��������e3�����F��v��n��ᚢKR�j c�u��.��N��\4�[g3 il��~U�8\�H�6��D�N��g�ԭ�BJ�~�M�6r�>��3U�����@==V\�����U��-��i>+�ޙ�ޢ�6��m�3���������� Z��BtJ�j�鸸�����&���@��r��5�ǾuX���h1ˀW#<6t�ҽ���,I�	ߎN�V�Pe�k��"$���+�u�"�<��� 3vH���kf��]u����@����|ͬ"���� V@��/�4pV?�$%?,}w͎��ny�:����SO��>ݸ��g�t�w�F�r�z�=r$�oN�*����
�?��HR�y�@�bH�Hd�|�O�
��T(C�dɒ(^�=�#D�2s�)O`ظ�-/i���OM7Ҋ1[돕֜Vv�G$r��n��G�ۜE� L��'53�WL+D��ލ'�����S� 98O�6녶�dJ�#��t��𒋟@^���;�1��-�<{������|³�	1�-�4�q�t��_ٜ���9�{Rp��T��mO~B���n҂vG�_�g�}jZ /�0X=R�,��T�c���m�!���Ҏ�`���L������)<��I݉��u���GL�1(f*1�(t�e;�"�{B���X����ޑk���3=��$?���>ӵ���F,��&��as�0���i��U��P�@�����6�.�<��ꪭ���d�L�$Yt破�
3��Zn�b�y�e�^x��[��D?���g6	��.f�9h��������{#m,nv�(�(@Y���ËΥH�%s���<��:��Xq�oW��o���o͔%�e7���"�R)?|�`�J"�l�ֹ�Vbq��Ş�U-3+��� zRr��R�gE�j�Y�>�X@ч��$���HE��-�q]��Q���!��NfE���5���ЬUV�;s�UKC�����!�d�c)e��o%�Įo!X>҅H*7��vW��oدm
N�����D8�-+�2��h%�F���]��m���2k$�v�4���\� I��Y���,ؖ���c�~���5T���γ�66��������w�Š���
⪃Q7Sxb��`0���>GҸ�)�AUh��'v���&<����X]W��6s������Z%T����a�Y��dS�̿��Y���R.�-�B��]R-3���(-��D`K��.\���ʈ���/��8�[���.?�E]�h�����]±#�Ċ�)�����۬Xr���c����M3 t0�6�S���(�;��_�G�>����X��M"��)|���d��>c��̛$L�si[��\3�M���"�������f)�����w������U��/y�U�fp������bJ��O�b;pu%/ww��4�|��b��mi+�0�)3��W���I`����	�H���B����Xh~P:x�2S��co��^l�^���QH�qT_gr(G 1cN���U��y���$��۱=y�S�a�R�$s/��i���rA�3O�s)xۜ{�7Ba6]<[�.�/�q�y�`f��}iE�L����ke��p���:��5M7J�mW![����z��
9� ���S�^����E	�V���1����լ4����0���Y���8SvZ���)_"4�$�Ci�kH�o�`b��Y��������'+���8(��f�Lw�C��K����ơm�U����9.�cG�I����9�}�����'�f�����DnrD���`0��јG�)i��PV�����)�񯤁ƫ=��Jt�����\Dˎ2������F[��@:�ELt:�A��÷fT��]w1����B�(��f���WN�2�m�Wݵ% ��yJHm����T��N��OE�����L�a�e]�S��{�UF��	4X����١R���1�|9�����]?�����.o��Q�w���%�	��6�n��|���Y�{ZL~G�_M,`��hc��J�:@�5�۵�)��Ih�&z�f�/�:b�XB�&�����^�?�9/)	ؕ�Sa���g�J��˿����E����!o-nI���Q�:X�r������}&�٢�wBegJ=�.��.`�nm  Ex1�����;G�n��\��R䯔�m�!�kx���O�af))���ȕ���-xbc ��~����$)���A $���:�Ţ*0ih��<Vb�!���2:���[����N�-�Mgr���=!XrD7��k'H���	Ҷ0 ֵ����%�=��?�\��G�oKk�|K�-a�ȺѴSʑr�5@��2x�MKΪ�l�����kq�UEQj�������C�����E�Y�)�Ɋ@�o��-؇R�� q�s�l�m�<�0\֥m~� ��s���&N�����Bs	J�������Ơ<��et��%`Dxߜ~��ۿn)Sk��OXL�
��������':fE5�Q���d͹ݩJT8�
k~K��+W%�H�B�����_Ʊy	��ccXeF������ܬ_��Gt�q���&�%n�3�ʟ>ߪֿ�� ?Yb�|����;��l!a�	���wȃ��4�m?OuC�3r^9��F��pB��J� #Sh�S'�h�y�����]�(��
��b���G��_F/�+x-��q�?�� �nPqU��$/��#���DZ$�P\q��Ě�)Wq�7zdr���鿟�?�e��++%B�D�Os�VPFpXc��w�/ւ�2DēcO1^RX}^���q����*����j+r������	jk
���aE8�w5X�L�7Hʩ�Aϩ�>�%��$�Nح�H��IhX/t�g���jZk�o��,4��~p���T��\1v�@fu�u@xmI5�83ˌ�	����_�b3m\���-��B�cD�j���� ���TB�S���P��H�~=% ���f�ˆ�C�{����wjN{�-�ɝR��94�}�e!	z�WG��A�R��/��p��G�)��(��N9%���_^��5��p _M��#N�o���j�?�~��/��R���򂘧4_�+����hBkU�7�x��/�/<A�����F�TWs@�Ҙ{�0�w�R#�%��&�]��` �D�+1i�:����2#%�Sr���K֐�Q�p��O�B��`��Z�5�>L��n���=�L���T�wĮ��s����ִ
����J�o��/��H���N�OZ�ଡ��;	9HW1P��]N�ko�B��} _V�  ��r��ķ�)�Lf^增�vK��m�z=�:��հ	;0m8�����2D0��\N1	N��u������D��_w�XR���h$��<+���}��?�]����P�ڃ;�Z����5s���R�x�8܃"m�oDk��Q �Ѱ��,��%"���.7/9��fp e�9�lL��!x���?���l|7�Y#/L%��b�}�E�*�Aゆ�:��do�9r��`���� �B���.MP��´&�$����>�� ����C���Qc_��\��x��0e8��;�?��CSA�Z��ng�A�k��jV]�=�of��Oڪ���=��}�ke��h���*01���l�p��`��~��MQ������ ��	֮u$\�'�(���&0f��<ݻ���]���2�S���W#Eu��_�w����G����.'o�)��� ~�/�^ocP�{d0衳�Z�7&M�����c�� ��EH��;����[";9�"��_�� `@T$�(k�X:=�XXye�ɻ�P�p�<?9\��c�P�9t��e�|T�t�P~&��z����,G7N�Y���B�9���G�U����@��F�'u�o �B�^�b��Y�2Z�Ѓ-���N�^j���~�x�,�������_���Od@�;�k�h>^\@+<�DQ��*?�Hџ8e~�4b��3��6���&�� �A]��%αN��[C�ؖ�_�n����×����t��D2<���"r#G�Y�s����K0���	��sV`ʒ#+v��b��@�����r�p��F��o� {	�g�d�+���$ELm�r+x'����	&<g�vq�ے۶���arӬELZl���u�o���a��w��[�P1sMy�WWbs�6e�x+]�Y����?�0A�f�+�v��u�	!Ѕ��c��'���k����g�Ԏ��vz�kj�]yc�Ɵ�-)4��5{�m�jN���J6A�3��s�K��^�co�x[fN>�-U�|��z������sl���NG���j�����/�9I�K�"Q�>;G?�x���������mt����)]�4p���'Ds��#<���tĩ.bl?:IKRGN4�5�D�+X�w��
c���jY�>5C_,�
��XTEi�~��_���2UxSI�7wu�J�Djs�_U���VB%��A>j�%H\* �7=��_~>ܺ��c����D�#w�akr�-�8�s���AY[��'6�h"��X:JU}�ܕ1~m�q�ؼ��'��Ӕ~G�d�����4��%�U+�yUK�W�1<2�t}z��_��.}�]4>��8L���j��RIw�G��9-:p�v{x� C|%�2|u�w>|�&�7�{��N�'F����镞��ƙ���/6�ibCQQ�R�^7��mcbm=*��q��:	�uI~[A�(5'VD����n ��A ��"e����ew��M�!\j=8l����KHx�>Ҷ��"��?7Q$o��EY�a�Q=je��=��{S(\Ʀ�Ø�5"��}�H"����k���<c�{�f���]J?�XhGX�%^�۽�ju1�,71d����}����Hj���ĀW�fh*�rŀ�<-��#��X�Pp�Ǿ�e��|՛��%et3���n�y>�f��m\����sj�&�����s���&�O_&E�,�����6�hnB[J��7��5�m��e�*C�-�JZh��+�K0:�C/���L���M{@&�6t;c�������~7�(�W�v;�����o���g����Xe@v2\b�%L�^��Qh��\A����0�vV��]+�i��wy�:G�Uz���������� �L�������K]A��[3��RAʃga����O�mIZ�V� f�X&��0ʾ.=iT�?���^쿪'�^?G��p�+�.��E�n�ES��Y\op�=��sNZ<%L��#�k�G��ZE�����!z�mH���^���d���&r�6�Q�Pց�}ܺF 9
W%u���` *�ߝ2TGL�s�wL�?yTK��k�V�큂@��Ԏ*5�6���4 �y���0�&�Q�k�<�2�������"�5�c=��-4O�3j83,�!t�_l�lk�%晿�5�FaGȳ[e���m���44��	O<��o�?Z���0�)?�t����v,�TU���r���?�$��yM[��)nÐ?�4�ZQ��&���;£�O�� �^�mEӞN�3)�z���i;2���ģYa�-�O7����W�[��Z"��7��m��]��EIի�G��Ԯu�}?�ޓX!]5�= ��Rm�/�t#�):�#1V�������~O>�ޤ�w�r�@��r�ǎ�$���1�!q��N��&r�i[3��vh�Y'���x�/Fq�\Uu�p&��5�a=CI��Ă�yuV�+�e�8�V+�,\JGNx|�9ZQ�P�Ȕ���YW&;J�J_/�$�~��?#aη@Odz�b�K�?~��R���S��
I�/��c�;u�����V6��Q �hj�pă"@��d~�B�c˜��������Bt�r�Tx���`S�1�T�@��Y9"lf+Ϩ|m�U�-���ٍ�t^�'�J��[�[ͼ�;%�
ǗU���ŏ�0t��{ᐡ�YHW-`�P���81�C��f���V=�����E�?�̠��Q�Ti̺b<e+�C*�?�Ь�r�I��Z��06 ?�'��⳨Z�Ʊ�~i��p,r�Yڽ&؛��zd T*�$�e��*�(������@F%tt=�!��5�n'h�g��ڊ��1 @��>]�0��%�R���k%��;������ ��rL$2�B]��gR�?�e`��
|_����NP`�ٝ���W��Y{o"9:p�$`  f�Ʀ9�G���s�@�p8��������S�+-' ���;4K"��(���	�7�!R���Ρ�������>��;�1��rȁ��{$j\�>��H�ׇ�!l�|���y�J�2���ל�5/U�0��U-}+���L�����i�u �~��CEk�/+�c)D�]V�>�kV�۟]�68ؐn�_�(�U�T�e��j���i�@�]��7N���L��u ������ g�3ja����'+��(����5�uT�CWN�Ǣ9/�zHv�1�u���q�p"�*jx�"w�����'�5�v{���!h�`������i�+5���MVi�>�g+�����V��ҡ�G��.���:�������Ȫ�Iڞ��!�Q&%�=wHN�C��jewJ��Q�?���1�v��"|�F�lO�m���|]�7���\�Or,��G�������i�06GY��b�J���N��ؒ|v��q ����,�{�^[�ec���Hj �Yy��(2��A��_[,9
@T���f�$� ��3@<>6����k�P��?�Z�Z��͕QR�����W4*���VE�_A��6m�k=�%���h�+΁�"8�Q�����įWN`��6!����	�\%��c�%�HξX�qRC�=?4d�U{��d\2��lb�Dؑ��rH*���z����8I��||�Q���ā��uN<+)UK-�;�!CwfdL�S;[�3��Eب���ީkJ��4ոq�/7H�<4�����	��z����� %mth
��������$�j�Y^����7nƶw�v�#`w���a]������[�s�\��W�����T�`��,B]��`������5��*�,�pdǻQ@��qz��}����^0��r� �#���)=��j]�| ���9�t�q@��>ԞIJFb3m�`| ����'��LM��o���H5��"�Qz�p^k�:"�s���vŔ��6��s��e9��"���ب���"���h� �yÚ)���sU�m��X������%(1��a�حx���:�a�;r��@$���Лy����K��Ws�m���P���`V!k���'�q.] !%�]�"��&��Re*݊���R&����hݐ�b�e�6���T�lC�`����_XT���o�ކ�� �t�g�`��d��D���2�d�/���Aڈ�wvk3m���j��em�hF��M�F䨼Ws"$���m��"0X�]�aW�@V�s�p�L3�,���L�����FtI���ʭւ�\�(fܯx�����>3��}!⤹��q=>��r'ܥˍcؽ�Pxq�0� ��N��y��/h��9t m#��t�]	����L�^��`��PQFW�wS���j�^�Y2Յ�Dn��m�'�'�8XA��6H�ʜx�)��:��ϖ}�`ˤ8yF:�x
![��=}뭦���C)������5�xj���7/_�dx#f���ˌdd�iXT|�e�MpM@��.ųx���o���v (�ڳ~|]>�k���D֯f+�O-&�Ƴ1P��j@D
�.�b�Q��0�D�d����4�|d�����0ީ!�����9-)�����	VPqJӁ��9��#�Q�a��1M�j�Z�	����3������5���/��C���0�Or��c�{�O��|��M�����[�#���k6�6<�49��.V�\�t��0� ,�	R�}��Y{�>�,�q�|0^��؋��m��\��ZPC=(��;�U8@�ƀ��4�e��#�N����30�?��d5�p1�E2������d$�}r��(�_��N���ԘO�b'���I��Q��ꈣ%aqP�i1!�����%ࡇ��cÂv�س�ǟu@�:��)�q&��`��A���5`�/8�ւB�>v�ז��_��r�S ��y�]��)��t��;+�Rt��!��~qm]&�k{o��>>�%�aa�d[���W2��5HZ��?ٲ �.u�KZu�����Y�G5�v���u�~�&�1�]wwx��Z��^�hhO�)�)zF�|	���!Tr�,���-���#��M���Q�t�r�����m�L�/��~�Y�=���#�破*�n1�H��XQ&C:��(=A��zj�Oh�#)���@ʄlQUdu0�k����L�:0p����<[#&͔����ɼ��d����`"����ʀ��kU���є���J�o;z[���zO0�����O�n�M��-v�I��]�����3�L�K�=�5��s}~�>Ɍ���,��l�.�⻫l�[�ؓWǋ�3wIܤ˚5��Y����|B�H���ˢ5&p�.�䟣�(�6��ܰ��^�^��8S�!�yM��gsE�������,X��7I�̠$������~�k��l���ܨ��Tf���>l���nQE��Fp��\�Xp�<U����Q8���H�9è���Gy�H�z��׌����5���(�n�� 6f�R��'l�kӅ�6w���R~<���3�.��-�gl��l�ּA����H]bL��8-�ކC�!������t�ӭ�$y{�;�Ã��,��\�)�K�z�[�QL�WѤ�6]�ݿ��Y�ѳ�V�A	���*�-:A��K��OC��w�JE��Vz��T,�ub����y������S��zKjGg%HkWW�DM��r_jA���꒥]�%@[8�}������A�A�-�s+]jˈ���2�j�L�A�	Z��`�m���� ���L^a{`��֗mw������O�L��6^}t�=�$�F�n��O r��2Ī9\4��В7��HI�jA�Q�&�==?������Y1���~^���*��ˉ�%ᇢt	��s_P��3��p>�\Ix�H�ϩ4���o��$	M�PKT�q2�4���PF��̡5���nV�C&��⇿���b����D�e�S^��MLЂ>�'v�v;��`�}��j	�xWL�	b���yvP�i�F�8��fUz,,��ȁ���-,����I4��"B}��PC�
�^]�r�� ��ؚÊ"�*.�7�}m�4�^9n���j%��C�+�.�9N�����°{���xG�'K��09v�,\���e��̊r&]�y_���It�m\$��0�8�Wי"�`�Ͼ"+�l��RY^¹���b@�E���%��o����'�`�Z�' *��R�I;�p��OR�e�;爿rdC��YD0�X�Ȓ��L�`�(P2���̏�b���@�p;�<�c��8�,fH�H	z[��Hg��.0�6�-������������؜+��Mt-�|�$E-���ȁ��^��=����Р@��d.ɲd�**�����+oz@z6E����Kei#G7�^��"lcQ� ΩԄP8�xz�D��nC�Uŋ�.[˝�t��4& ɛuq�<���]l*u4b�n��F�qڤ���A�؁Na���Nb�0r����k�`�ʨ���6K�@�X�eW�O���	~l�X����^�X�75)H�N��v�{fR5�iu~ϖ,N�]��g�C�ߤ	�k޼��[5Q���\����� "k)n�88��Fe��1y���l]��3��u�1P����rH���*+R�k6�� Y��5����%�љKO��m*��5�h�\�c���)d�H�9����	R��b	Ȟ�<�.-���B�O0� �z$Ͱ��Pa噠i:��CN$R�տt����r1��31r*�h?(�}W+�fL6�����|�]�^�``{�ܙ�#�'��ط&�'3E���vV�?;�̯jN%��}�ބF[���)+[�aHfp(�H��z�u�	W��Ȇ�gd̎�WD�� }�p�����1hR9��a��>>�ќw8F8���������J�[�l=�������O���c��>v�h�H�ǆp�Be�3�s�h�I��#0����ߔxf���I�b�D�K�P��l�T�:��Y�冠Y�JQ�
%ߣ�kU����~�ds/;!HϜJ?�G&��������5��(Q�{���"[g��AA�b5�+*2j��.x0�k��7;HWf �RNy�l�o�h�у�v�k� c 5}Aw�/��y�6��%j3{p�
{�*R[	�?�Z �=�h�8��6���x4/������-�[e�Fr>��_�#�aK��+��O���
i>!"'��7~��ۥяjx��!���w��������ڦ�t	�C���Vޏ�%"YjI2d�w�V}�d ���]�:�C�!vϴ��3��O��W'<��4�-��-������A�-�{���V��A��Q�;�#lJ�>g�����xr[�R���u���>(*y�zi4g.�p�?V�`����.N�u��d���!�󲯚�m�۞�q)V�e=*���H|��_�l�nm4�MR��7��1���N�e�U�(ҋ��6�|f�m�Lo2A�cc����U���d�H+A(���µ��|��n�I�._��� ��'��Qf�^'�d��'� ��3���\`u����~�@�4e�$�@���(����o��fG��TA���e�����\H˃l
�3������ۃJN}î;��[�o�g�PV�B;�h}�%wn.^�(�[���2�3���hxqD=�7?B�
nS�RI�z`��q8x�����PIcu7b�a�i�'��(�_�L���pt`�~�s���!�$<EE`?��Vk����ĄE�S�c�z)��b�W}8?���)�v+;����@h��q���q��e�Sݷ�*n��t�6!jo��p������F �5ߜ��1P޵��>��:����1OZ�#V~���e�{,=�B ;�f�-�uR�P�� �z��v��A$ى[�	֒Ԫ�=c6�JF>��5�L� 3,"�I���'b�Q�|�ꖵ�^[���$$�>�!`M������9=m���A��kN�\�G���"�m�]yO����獿H�ƳqqՒ�L�X#Ny�^�猁Pvc��n�dA�G����U|��N:I����Xv�s,tg���^���;��
sM���~
w��&���ʦ��ۮfv��5�U����E��#�7�֙��۞�g$èk�F��BY��Q�bJ`k:I}�JWn�	m��)�5��b!�d�x��I;W9x<��_��[��ٖr2+c��g�F0�ܒj7�N3��yu �|�8RC����G�ˮ�������p�O<U���S�D��b�}�\�$E	V���uLz�ՑZ3Y��)*�������:��!�K���&�-93S��kL[ñdq��焫|(�!n
K\D�r�;TO���\ǂU��M��|�ʬ����!�h�o�~;j+�C�ZȮ��,Qs_?�Q��|��)��^!�{9�����1W=>�A���aL����Gg�ˉe�4�'-�x�\�B騮�_j���U{,���L��`BL&�0�^(��VBC�
�.]6�z��1�*��l��_W�)Kt�8v#v._�<z7��f��y*�M�#��t��^��s6�`���9r��ّ %�05�}Ul>�y�)�K��.>�Tʇ�2ط�_]4u��z�����2J1�A�:3��)� ������%����O�����G,��*��1̆�F��Zy/�I/�S7j�/��3�.���o��&�n�_w��v����I�|�I�O�B��B�O��ئ1{[������Ǝ,Tǁ�>�c��A	��2�bJ�Zw�r�#n�)_��~D��x2�^������eFDY�HܪF��U[��O[��rI�U��&8�q�Qs�`�¼[oJot��R'�Wt$��i���c���e���h�@Z���/#��<�D�������dN~���l����U7��������.k
�s�%o��Hƣȧ�$�dD�D+�Zi�R�0�=<0 Y�W��S�!��3�2$��.&�xy4�jT8ݪ^���o��%�W ���'r�?`N�ԕ��	 '�q�|�Ť-�rcQ�?MG���#Xd��Oxo�rפNV��R��F�W�d2ƫw���v�j"Kp|?~����X9�����»�Y��,��t�&|rMg���	&�TM�Dr�2���7o�LyM���v� n��ֱ�:<��
i{� ���8R����UV�l���JENu0�of�e!>S�J��!o6ch\�S`����B��^�z��s�1�U=7EL��a�C1Vf�ݍsf7��V��~"�^V�7�:��͸�^�-�yV�>C�������A��Y��F�|c����w��2��W*Q'$�U�*n2�Xޘzr�ڣT�*|��fI������s�}�S�@U���;��	���D�c��W�:���P}���Eي��vk���.e������q,OE�DP,�uk.�d��[ⷉlt:�Z"IZƌ3@�7��Fn��t�ܬV���<^�*uW}[�r��Vf��Z	o�':'&����ź O��M�6l!��N��E���5�h+�~�dR���nL�X
%æ�A&�/�X�;$P��s�(z��A����`��fׂd�����t�A��A�bVZJ�n�R��Q3yL�#;13���S��'
��l���|�­[ �'
5�f�n��5���Ei��T�ꦰs�`H�G�����/��4O���N��
��'Ve�3�i֫��Yv��nq�~ڠ��쁝W��ѕBY3�0�Os?��������0���IW��vݺ7niaŠ��Iዪ~˅x� y�l���#iʾ���{i�?h���XP�B����L���T�� Ke�`���1T� �F�Y�$�ưFw��7{��D��S����N�w�G[�s� ���g�"1ظ��acY�zWף�_��I�*$R���H����^�'�>�Y����g���|K��	BK�v�#�� fH+�&��t�Ȳ,m(*�ͥxQ>dh���c��S�w��ٸ�ߥ��l�[.{O�3Gm�>N<�ƙ�"m��\��GӮ9o�3h���{m�6�������?�x)E�����Z��ڞ��G���N����j ɇȎ濙���\�Pcg�Uc�.7a�7�
�`?�����j˙�|�����Ў�+�����#�u+!Gxb[��2���J�4�s`����X��`�8c��/N�a�l�\��oS�A��AdK�P�k8��;����B%�VG��NM:��:.�>�h~����0$l�C� ��k`�cpf�G��o����!}~��J�joc�S'��RZ<'O�0:N�1�o~�����ca��~�h!g\'��-� �Khz�Դ���΅�.�����0�Pø��kV���(��9}�^E�.��tp�x�����~�狱����P��y'3-��_�Zz!9o��A�_�}���x��"��!��Ϡ�HF�K�����@�xE)}�������!�}P����T�kI�q١S�;)�R��a�G��]=��%�aaa)(�'�n����ozΊ\�En5��Z3-vYF=َ�����^���!Z�M����wf��j1+c��i+��0���:�rF�9K,+Iw��v�c��ㆬ��9L}�B�݇��<�=*��=(��1�\7~�e!׆jo�{��%���c=��k\�����FI �9U�m���%s��pO|$�A������d � ^���T�-�.��<��C�T>�+� �,#
}G	�䨡�7Pi�wG��{�m�.��K�L�k���!̅m����04�b]�� ;)�;������z��r�ȝ�s]�����N��J(��cV���#(�Q�R)4�R 7�@6T8���+��8����Q�#� Qlì>�	ڻ���	���x(����kT���3>�^�"�,S��tp5)����{�J�Qkg�6��2��L�=��|���o�]��h/��$_X�#^�h�V&�����(�����;s�v�C�l��-F�z�^4�1a�R�).EUT��%$��V�$I+#:�q'W�o͢tsn�[����e#]x�d��o�aP��W���`U�`̫o5f�5t���9ӵ�4�v f��\l�~I�yo��ӣ?R����bUx��ɂe�0k�i`
�<��u�p q*r�K��%���"�D��vl������������W:�n�Z1�z7=H���|)�daaH���g��PV�uh*��]�b�`�� tm1zg2��OoO}X�59z��&����Lr�m]*]���yV��ހ�5�,�{���ٻz/v����Y^��09TyD�x�7e4S����k�?0�De�Q��u�wv�w��/2�i�˨��N����"�������d��g!IN˳\�`u=;�~�������x=I`o��gk�h��_�}���1p�H]9�p���]�8Fg�䶱I�k<�O��6I���;�^V&���NR|��U�Vj�f�iYN�r� �W@��V���}�~�M��ͤv&	��uD�-��c �V�m��	J��G��Nԓ�/�_MD�~/uI���Q�$�A֍�����eթ�2���p:--��T�Z��	l^/�2��oN	�"�f�e�Ø>q'�����:��)?���i��ت�V}���_1g��U��}�y����8�yq�+]�lp"�f�h��uQ=��jct�+uLlRŞڪ�����e�M[����W�-Q���+\����j	�4�]��cpl&`����kpQD�!�[`K���9�"c����7>�v���A�;�M�j�#����9V��+�sw�>6��&t�g���"3���4��h��eYqr�Z�9@�o�����C4��`l�@�{���,���j�aG������쿱��	b�,�y0Y�w|������"V���{�u�e���9�8��i_oH�˦XWB8���{��|�����C�2��yH7�S|���|������~\�+�B�)P�� ��|�� ��'�5VlTj�/ѹ�Ə*�@S#.�Q�S�,��7���<3c�5S[��s��K`�&He�i]�����d�׽
}琷Pj/� �ҴNȹ1�Ү!D�.w:J�H���q��VM;�1M�����@��a���B@Q�'�C��s�����g����[C14��1���k�ˏ�h��D�R �#EVO��ڇXmL&���SР]/U�!��Y6�N��|�)��{���Z�����W֏���͡�`
)���UkNe1�.�A}J`��"�|	�)���{ V*�]�;,3���k�q&f�w奘��1�Q�7�۬&�^�s/�w�[6���,9��hj����]|ߊ���;" ���اޕx��F��(o�#VD��s��u���Z����H�M��,S��"e��v}���$��°�U<���!-�Y�A�{������c�O���[�gcwܓ�s�Y5���&�qx)-��̅��`��in[v$���xD��}��?5p�@!��[�*����˺h���+� ��!q�g�D]gɧ���i���\JV�����5蚚��Βf��mա�y<�即M!9����$k�nE�3 k�q7M��D0��l2V��/������đH���'o�丣��EeB�5��{�1�����yH�,T�f�@.+n>�����u�b��v�&u��R4ݱ�)�Xـ���d��Xeԩ����w�rNm+D[�s9/8�+\һ(�	�f��)���9�ӖGJ�B�lhM�NC�H���8�����&C���\��[�l`1���km@ѫ��Pq��U��Ѩ��ܑ>{��I�d�Ж�UQ�����`��s�-�z)L&�_W����@J�#��D�S�� �Ā�|�y�ף����?S��� ��Τ�%yCb��I�����|lR�1����Es*�I8��r֎M`����>F�����<o�o���&[��b0�ɓ�GϾ�CPZ��#�Q	����E2M�7���w.#'������}RcP�� p���V�K-h��h�M��A������ހ?���J��6��T՞�r�9��x�u��f��L�z�-�R�H���v��^�Ѻ5�\ǰ�S΋��u����;X�G�m�=���nf��S���)��B��Р������sw�*��_k�g���z����X̌eno�� +D��$j��\²��4Ie��;�N)�_$�!��I�+j�A��tG�zBs��A�2Ծv�� U8i1mc��e��$
d�Xu?B��B��#�H
oǐIh�~�;^z��D��l.��p�V�3��������/��VU��p�&g��� ��#���b�v^+"�M�v�Tj�v#P7�N�/YI��Ľ���!�Y���Z�y��j�%i߄:u���2VS�g�W_��˖1(9ǂWd��t��Pô>ל����|d�"ό��IzJ=}Y �k3���^@�X�鰓��2��֪9�9�4�2\8��4�@s�:@=����f�%�j�"���m�dT���tT�u5�o$�m=0e(��3�ը�;�`�˼v�j��Ȑ�2�=Q5.��r�?�B�#�ad`_#��&B��OZ����6C��T-�y<�3�-���A�n��rZ����70�ёa��&�HV貧vX�~s&fx!L <Ɣ�/o��/C��;��0��&�4a����5��9��/�T��t:��X�̊��/~e���'�+d��M�\��T/�3�&���^R�)#a?p�e�Q��x�����[���h�}Ka����mu@����{�~9'�-��f"�rOF	�������Z�@m�Yl�JWW��1������1�ʗW_�����
���,���
�O���)"��H�B*��X&t�(��Ƀsrr�wĎ��.�����l����.q9�)G��)'�{:J�(QpuUOo339��i�H�Ĥ��U��v���3ztJ+C����jV������V����αW��v���p�p�]*L������[��h
neP��R.2k[��x1|�C[�i� ���^���	�hgGӅYTbKbMAm����1��_̎6��Y�q7gUm�]��:haꊑ@x6��)����F)�+���^?d�F�r/i�X��X`_'ƅt^c�҅�:������)"OQh\��B��p�r�!�N�z ��wtb��W�k	�D�i��әӏ7r鈳k�L:�.�V�.K뉯H8�߰
�?.��"�9�k`�J}�S@�$cɒ�7ߠQ/T��R9e�V=���O�j 2!I�u�/	P�����.Ğ��W�V�"�oG|F���p���x����WN�
H�v����%�d+S��k:���j�5�Ksqe����YDp�r�w�w�a����1�R\-L#���BZ)�0���O1�%�DzV���	�P�#�����t@��2ʀ�S¶מ����.�P�Y���zd����5P������A��l9���r}0�l���*��*�u>-��嵵ܙe�
{�����l
�K�.�V�k�٥]����@�T���7�مI�����*޽.˂Q�Nkr��eF���sFq>|�>�����,�Np��jL��ʔ�1uO����߷�u������7�p���*̈́�-�⷇d ]�o�>eGB�
��d�2+pí��B���/G�!�?���k�?��;�SFdq�P�jv���F|�ZC�vj,���uf5$��_,� k���2μ�����bj�ydO�1;���1��U0�0U�{��}�puw��t�O�!2[���7��~	��H�.Y�eF�	{F��=����[��i	@����/��H<F�������1�<�2���Z���]��A1v��{w�Ã�j�]�E�$������ �g�/�w�\7�#|����6��R*���ӦL9� K�#p?��%8ì����#��}Rq���o2��痒�@������8�j}�m�?jAkKyb�j+@Y��Bx���M�&��6���T��>C+�E"��"�x�ۏ7�;c*��Ƅ�`m�x���^�6�Z�Mn�6,9�e!�RK-N���� 섟���|�������W��γ�a*֊����C֗��ih�z�'��L��$]�#e���?k�E�Nx������[9��==�������B�U(�j_��uJ���% ��7h�V��z��+�X{�,�/�wᰱ��0:Ͳ_��l�h���(�Me`��v�b�b(b�v���`*�(�ٯ�x���S���
fNU"3
 ���#afݸȴct����|�e�r왙Z���E�q�iGY�g?�Q`�	?��KdPq����׃o���i"T��`KN�m�5k��`�<�m&}.��i���?���=ȳ���w>b�]MQ1τ/Q\�?�o��xX�ь���踋��0�ɩ:tшC�ߏ�����Z�04�Ľ�>b����o4� e�\_�<R�Ur$��I��*ܑ�ҥ��t������9����4;��q4<�|��l����cM�E��� &��������J��1žw��G��h��zڴO�-��
%��T�~(xW�ު�}�|��>@��A&��R$/B/'YuK8�s�{5�u���qbJ����A�}��?c�>�]?���"�2�#)�\�\��3�B�8��.�&�q�kf���&k+ܳ�� �� ���-����\Pq�2CA�b�x�2T+0Ey,)%Z�ʥ���+����;�i
p��/�`��v��x�~��M�왱�O�p闠y�Z��>$H�1,1�$��; �.�P���:DF��Vp�>��+���?m$����h�u�%��	gm#\��$�Z����J����?��1�{��H�����y::>ɼ�8j�(��Q/t����m?hK^����_ ��v��*�@;/r+��Zg��!I�2{<@& :7|~1_^Ef����
�<>��ٓ���i�=x��BJ@��2��܋���1[��~�Z��Q0����7�@"�.?�H��6��žzuQ�r��1\�ò��e��>q��*�g�������Q_�_ok����o1� �s�ݢ����Ĵ@j?^7?�|ɔ���˘W�Ƞ��v��4M.2{ݕ�Y��>�x:ͽ[�]L~"p�=�[
�B��䴺���s��Z���`곸47���е9 �*��٢`fS��@_��zט�6�����Ai̳�����de)L�6����K�F����V���P���=���"���MҊ�ܕ��	�H/���r��s���^[-���	��}sf�Ղ%���4����.Y����&��sG�C�|��G�����)^(�J����-&Ӵ�յ�ҭ�9�a�bG���c#�*���I'��l�*�� L�U��A��LPP*`i�ȸ��@"�fl��Zv�u1��閒/�V}%16���R�°?;ߘ��4��E�2lF�!yYI�0�C~�4����U��!)OD�C!�]�(�� ^"D|��_f���U�A>8D	k;έ֭���F�� ����ă+0��:�/G'|EBUh}��?%V2�y������h9}���<y~���_����GO���!ȨE�O��C���#�$��5���3�~(,�А7߈mǹ�4��zz� ��R��6�߮�q�3��jJ�-!��� '���a>������!h��!s�^��<����-���Vؘ����o����Qs�ܷg�+�	(�/kw���#�` �j���lw�'Ɗ���[��'��zpS$a;Ǎ����7_a���ΐ.���Nv�\*����9��D>d�xƠ���jF���HO�����~l�zܡ��6���L?9^?>�Pd"ڐ����<VW�:����ۇ�cA?�\���1�������)�W��e	�ϣ�Lk��8<NX��b��o�ۓ����g�	w� !�������锣��e�����gc\*�Hce5�BKx��PL�ﲿ;F�$�;ϊ�c�i�}���Ց*��%�=L���I��YRQ���sdݣ5���.�G(-��ݚ����[.2J��(���[e���;g8A��͛����T���~��k��+A+�����`�ķ#��Y�B�yO�/��]�1�`��;�+���������7�;$��9�o:��EZ�}�
����D0����]��i�E@�)@Qb��0�x*�ÿ�s!�Z�m�����E��;(]Ew�ù���"#��И�����������GC;&�8:���e�L���V2�i.>�a��0'~Z3[]Ct��iPs���c9~���~^�%�$�6'3�캀83�!LR������Y��|(�Xi�Pk�=� �ݮ���SE��=$=��[���&�h��c���8��A��[��A���#�@Qe3�lY����.�L��Fh�;�^��⟐kk�W-����&Z�A�/ΐ�/TG�鉐�n�<���FL뽮�"E���R������Ą��0��c}�p�������	:�X�6Zy�jps��1H$]�z�$y������F(�&0��?HGҤ��t�_����ɧ�zS��$u�
Z;L�-�I�xP�K����|�=9�6�~V��0��D���F�Y�zlw⟞�=���-��<�=5��Z�_��2w�'i=UR�_N���Oө*���gM�օ{Ĭ����_���>�81���tx;b���^h�����ħ6,�P���`�2b�	�cm��t��� �z/b�k`�U�� Ʃ��]��ǰ��Z�0��^93S�yX���K@D��Z�Z �}rQM��4��]Y�1���Y��f����V��Yk�S�:�jZ��!�Q��j�#@h�]�??$��([����;j�V���k�)hPA�-mX�s܅�Nl����r��*�P�ݲ�=��D� ��#4�n+:8�N9 �$,��}���	�/i���R��Z7?U�n)�V�A����楞���S�a�H�����-���邓���ߥ�,g��e�V\��XBx��J�}��;=KJ�3�,t�|1K�I#���}���l��v�l��O?i���l 0��6'�����ځ��3bfAL�%i��w�s��G�F���w-1!�A�9����=H~�#�*�8��Wl\��&R(��%�����$ٸEe��s�0jw<���j^-�W(
���w�?��
iT�4{\r�Zmׂ�!�.^e|勜�װ��2ƈ���Y���+Eݳc��F��]ڮf�qx`���괤M�-�(�[sWGpQtp�2,�A!@0��қ�w�a������T�{��
�uB�3�,�[p_���Æ츧!�r�XQ-cf�{�'N�2�ݗ�8i��{>+m,5kȬ�w�I9F6}���o��\���x{�*�=x$�,�#��io ���ua�S;�j��C6I�f�j^���9,��Jn��}�$"y�r/W�Ժ6�|�!���,.�F>�?���bߝvOw��At�VF����,Qv[����>�(Q4����h>���VJ(k~��O��p��:|Ua�;$���X3�G�V��tR��tr�M�&�m��t&r�b����Xz)���*�Py��8韔P��
���X��riS�ܸ+�l>�q���݂;N}��;6�ABU�Nݭ�'6u�� 	Ŝ��/�FxH���c<z�ŋsD��z(���b�2��\U��i0�0+�c9�!��&(���n�8�J:ʁ�қ���՜:�m�*��?S��R�|X�uʩ(��U?�8�,v�:%����y.��z��y�&	��B�1� j.��E�io�aXBH5JP�R�78��S,lZîN�����σ��\�Hn��m��y��IrVe��?��}��[&+�	��tA{��� �(p�����%��U��)"IOPҝ���v<��d��5�\e䲌�I��B N�%��T�U�M�)R�#ɫ[����K%K�:'ʼ�^�]Y����VmD.Qz%�MfwG�Ȉ�e�=<�P���l���Z�+�Z�qU�4�c t]�cNdV�^����j��&A��g�Lom�	�q�k#�����ö�ĊH{Q�����"ͳҙ������T�ϭ��[�"/�\Ƣ�ϧ��s�Һ����.��Vn4���-����̂�U|����+���]ݛ��{�h�Z�̱�3z��Ok�_Oi#e!K�9Q����`!��5V��~$���6{T�}�3�+*NAQ�P��m��Rr�:���|��,�LVl� �B>��d�#�[v(��挴��(�ٷuOLJ��cx1a;��ͤߧ�a�pj�5��A��hOw��.j�<gE^��YB �\t�����a1�c���H�XL:8C�Y�!(�������7`�n�:���u�0SSdt�X�c��,*�ǒ�����c�}I�
�t<�J�@�-n�z}~��;Sʽ̈�Pt-7sưqdU����dI��U-Qx��"�H:�]�쑜�ypuo�ΰk%��61l��ӕ:-{�'ḠK�I��f.X�>s�|j�ɺq�>h%��R�SG%w��n��~�[��.mL��g��Q�>փ�YMc]Md��q�C����=��~{��1�=�筕���_`���D����Pȩ�OSf�'�q���4��+D������zj0Yr�7��_d���G[�=��ò���f�m\Ƚa�3��SG�n��T�*��G|C�9�f�w���9~a��o����^�U�� � <��J�i�A���h�D��Q��}�����蟚>�i�J�i*���GP�����U��bn��1�ص�]�����`�o��͖�ݳ��!3�����|��U\�5͖+X���e�{|{5gP��&rڭ*�tFW5�.ɒ4�aѧ����mWBk�2�����˃�ɵ��xt��h�Ǻ���jA������^��ك�"�PE��f�WT@����,��O [%P�F��[^�Wj~�ί��Ǉ�v��xi���9�Kʊ{��ʸ1�����\W^�����y���{�H[��13e�\mv����'�c����Jӣ�a�n�nӵ�۝�����U�TafR�ޯ�/��yy�6�v��hl��nS%�b㓴�O�sp`_lx��iG�"B��Z��B��9��wXȨC���'�{�K��a�Yꨧ��[iO��hn3�h��J��<�c�,����;��<H���+0��{d�]�h���=C\	O{}�{����*d_�="�˚�V���Ly�A���s	�~V��hv�w�7h\��q!d��~9���O�ƃ��rW���f������ ���լN�~ �|����b��Q��Y,B葧��u�Cs��k�.��6 ?&��^�{�p�]!8�>�� �T�:+'/݂Y������7�]����RfCG�di���h���ѐ���^�&D��(� ^�q�K��G-�s���8����L5J~`�k�mM�1[@)�qÚ
����;��P���MIb	l @E��+C+e��Ig���c���#/��8�ר;���^V_ ��ǒ������o�2u�߽L0���#9��m�Pb�Vl�)=�e�t*�{�O��li4{���c���Fǒ�Iow14�h��*�hפ��V)f>x��
r�\4*fu&m>���ޠ����X�3f��$TDJ��cKc�����ۏ���NQ^>��z�έ�>�I�w�ī�A+�i���Y��}���A����G;�&\���z?~^u��i��0@�nu���IQ�,���b;i@P���������]mAY*,�b+�уŅ�s�l ���U�M���X^5?96 �3�F�J�~D�� ��7yk#�\#��;�]O1�$��Ǯ���
}��gW���t��YL�AX���#�7p�@��54@\�����C�PYD۾8
ZE�-�Ƃ�FM�\�I;���'��>�Z�t�O�\�
����#�ZK2�^O��QJ��&���}�]Ş@�s���)ŉ1�x�1��;䅚 ��z t��+ܙ�ׁ֦.KI��~^?�l��?A'aƟQ�Ў5��{��d�:+Z���M�G�~~ӘzYA��G���r)Q�T��G�V�4�����0O{���W��:�;��R�w���6��dh��� ������wj��+U�[�]8��oʍ#���"&�~�{��\�B�Ą����ګ��Ɯ±;P#'+����Ȕ��0�!@����A�N�� #�6^b�M�!{M_��K,��~��Cq^{�M@g7E�a�y�̍���U�W�r߰>���,�O�zuy�dv���hW\4���,¹>�@�h׶g�����|��v/B����n�T(+|*�o8�r�k2�-+��wi~�,Ta�u���nxs6�
��&����)چ b�*˯YA9+b|i�e�oB� 4��ǌ���^��~�<��r��j�ʼ`��R�a3�X���h���u����XS���N��~Ē���j�B���L�J��I�-X({P�U_��ct�5"��j�S����|�I�B"q�3�<-���+4�׈cN$ -_�~�5I�����P�ot�Ʃ�N����k��e�fn[b%Y��{����Ȃ��t�*���%mĸ��1.e�RaF�斜�8]�l�-"W1Ѩ��)l;Z�$ڏ7��0�����*��(�,�x��(\m9�t�CSQQ�l�� 4+���z�4+�����OcP�����:�����w�v]K�}J݄��.�3�-���u��|%~��l������=l��^�4e�	K[���j�jqe`H�ȯ�k+��Z�Ĵ��}ԯ��a�rh+�h;)�:|ӛ>���n]ѸsҽT�4����*�||�V&�^rõ��6�rހ�J�m ���d84PICZL�+��=�<<��=>�Z�]����SP�R�;� �K�b����ywH���U��xB�eɭHh �`�c	��8�s,��5s7\�
�(bU�Ng,�]���I��_��3��j���x(��V�ɟ�2M�D�C��&	I�f�y�2���ۿv^��&�$|ؽ$+q�/��E�l�<�5"GYC�ݘ�/�((N�}��DM&F--'��s�A|;r���K0����.f�@��'G_6��������1>���V�[&�A��+�Wql�l ��1�aH���`�O�d=w�J|���]��d�"����r?���_Z%u\to��)_Q�j3�a<���
��iEkI�Y^�4��v��1�D ^
���E�7�#l���- e �+x��� �A,%��AB�y�����H䯔2M}5�gΑ��$���� Z �WRX>�6v��1���z�ik_�����-�wKg�5w
ܻ�n?qU�� 4�>�������ڪ�	���U�_�_��ܲo� cjuCj4�f��2�Y��̚���b�		�͞�����O�,в�I��������)�8{�k�e1�Z�����%�zW�#�q��ݝ�<g�\��P۔�I�g7�9 �~ �iX�瞦������>��)$��CvA��!|)L�-�A5���X�^fY iSANAc;b��ܣ^Τ�^���)%���Յ������y�u �ڮ�䎘�6$;�E@.oo�M�JΔ���^t���ŹQ�c�\�G-���!�)6ج�J���RV�ʑ8�ijϺ+ǧ)��W��;����k�h]N�ȾV��� s�(�!���3K�ь��b\ȳ��t�L��׵�V>�C��%;{�1>b�r��w�P�����,y��xp�"�ݓOE�۲��慀��!ȱ��
Lj�]���J���;S���R�w�z��>L����]��Ͻ��$!�s�	##7Of�i~mWF1۬+�͝�za�J�p�y]7F�3b3�9��2C����s�>�4u{�f�f�q9(�V�5�[u�3��<��Ə���6���GQM��<���;��]��Q�f����sOf87,��)]t.S�#�H�zF�RV$X�`���#%nҠ��� ����<O�)���F�S�R�r��HlOc�<(��k�x��ǖ�5�w��c��,J����(˪��R��G���N |;�P��iR���[{��4��m������-y���M�NN2�[m�̐pE���l�<��jĴss*x@EH�h���q0Օ=�[��@��u���n�B:�,e� D��d�1�݄O�w(��#�9�%@��M�iwJ�]H/~��1K��ѠY�H�c}���=^��з�l]B�:�9��uL���ƃ���H��v��/���p+��bC7�<<m�๼;�x��6�w��W)��k8Cs� ͵B6nk�Prb.U�c���h�N��񷶟pUNO�CL9���ZyD�.�9�n�s�ߞ4��=P���9*�)�K�{Z��$���W�%�	]�����(U��%O�j)�ַ7)^�փ��f�ΕV�%H˯�(�J�ӕ���l����)�=��ߩ��x��l��s�t��K�gZ��<S��c-�L�PFW��xgw�%�U1��A�{&�YeGh{ڊ7�kc�Z�NJ����og~3 ���;#v���M��atu �������A�je���+(9v~��	n]Uz��V��C�X�x!�V�J���p8�|�� �j/��/+C^�R�~������uc1���X�.���6�#Ȩ�5�|���9$���w�i�o����]R72����q�^��ͩ�� �����TB��2�s:�ɛ8��΂t[sSy�WylԹI�}ֿ����,����#5R�<:7�q7]�������j�OP�0�E��p���
���Q���Z���UXI�ƴ2x��I/���`>�nُ�Z���n�B����| ;7�-�lH*��{�=�������Lv�)�Y�2�M�^�䴸�	�r��Ɠ�DENF�x(�z=pV��u��� ӷ���l�8]8jr�k���=0���x����p��,�1ǻ�?����?��;m�Ol4�Ӣ]��g?!r/av*�P��#�� �Z,��	��k��@.��8��_�����rA2�s8�����"UA���,=� t�tn��a/���	�v�.{�r�|XD����.`ފ�p��=��wt��	
 �OJ�n������aܬk�(?�n�9y��1��Ѥ�h�#?��7�B��zM�=��;��,W��l�ԭ(�3O�&5���6��sݤ�;t��Yŉ�j!�cL�-�{?���q�3�y��m�����҂b�A��+����W�T��D����J�֣���>�DL�p�l�K�8%!Ⱦ��q�		pa��3����ᴢ���jHmܓ�+�Gͱø�Z��'/+Qq��-�'ɧfNԩZ����e��@�إtѸ�e2/+�ȥ��iמ^_��zA��59jnR�ٰ!�Z��.�KN�>f)l&��"YyP���
i;��31�	��[��~�^�1�71ءG����h�י4ZF�YX�|��٬XS�M{U����NyԀ�����&бX!�	D/�p��v[Vir�d��Ț~�O�� )�q��g��Ae$`j��Lf�n�<�^�}���a�I�K),��������P̬���op�<��-�!2��b͘�)V��ۈ��g �S��ky�"bk�-�B.�A7%}K�6��M��]��He��� 4��]2��F*c��5���񛷏{D����"�J�E�tП\e�ِ×3��u���X���K�S��m�	�}\듀�uM�R��!�1�Y��Z�2@\�u
ˡ�� j�������n�L��Չ��o_t��4 ��\��'29"P�Бq���ۧ�i`�gU�/|�ŧ��8*�7! ڙ��2�Gk���?3ԩA|ͦ��Q�x{�l �z��-,-��L�A�u�U-�F��h)��q��r���j"U!G�dd����+�#�@ҁ�X��ײc~�}nawJ3q����rg}��s˱��ʋ�r��,Zb§�Q�^��Ϩ).5f�}N����d�pE,���y�WI<�aAX��r��#�����2�^��_�.����<�4��j9\.;.�G�� ey�s?�U\�}���7��k�#~���������N �u�zP�I�u"g��1T�Uc�$A�Rp���������c
������L�*f�
u(�m�����T� sNe^?h��E��N�g3�Bs��W��ɚ�pɌm:�,��B	�A�-aF�r�cq�l��,����c�,PK o��	�J7Lp��P�P^�
�Q��\B�PZ�pƆ�9�����P���X��vͯ¯rqz����H�^�$��R�)B=�ܺ�)]sT��IV�����u�ۓ�_T	��XeD�2�o+���/�G-��)�{q=�n�nS���l��������]��/���0��ΔԵ�MH��S���$�/�� r1��ۇ����9X2���O!j��F�6�J�̋ e�CT+d���s�$�Bp��>9��R*�j�;p��:x��2�p��fq}+"�]ڌڸ�ʹ���祧�Hg��Z���~�TZ$���� �s�K��/�te�kP�J��ki[�ڿ���ml@� w��LX0�
F����X`p�P�$�|W�0�.֫6�+�� ��K3U�CF{ȋ9�)�sL�:�� ��ĺ�I�9�{l��t���3d�s�b#im���xx�R��Ʋ�J���֦�ZV���C̶�W{M����	�Sw'q&�.=����V�y��F�HG,0����==���V����y3�^W�;�_����NM��[ ������ZE 
�vA#�K���52"�e��Ϡ�;M������(hĪ'�\��0/�5�1��Ϝ����\�UdZp:H��]�(.��W�*��sU�,\չj�q�Uac�6B�>�H>���K�ίw�:�]s��:�I�_�ul�JІH�񴄐���p��5�	'ͅ��6��)r������Y����˝����v-��S�bmW�Ee��qJr����ml��ڡ@m�P����^+C��'�tjh����Cw6�&S���>��<9>�I]���t�gw9����>���;c��US��{�v����luaĕ�%FR�`MW"�'�I���hF�$ �@���u�(!�?��Ċd�h��~�A��P]�iЊ�ʍ �v�<}P� #tg�ɋ�\��a��n�s�Jy��r��2�y�����38� �&�3�9ffU��U�[�t���B�	�`��m���K^e�
T�?bn�c$X2U��>����Ϝ;����$� ����Y�9P�;/E>��:�!yw�!%4�krl@M)�m��Q�Pf4esWVj<�R<P��2Ht�_}Y�i�3P�%�{q3�3|{,u,HVAG�,;b����&�;=Дg�,p3M����AO
��p��C[pI/�m����Dg��Z�Ĵl�0T��yJ�8�"?[Q0���s��Mx��<x�\nP |�m�dW6�)�bm��!��=�
]�ybN�O1�i��Tv��Rh8�0Yꨰ\�':.M�iX���!�wP�r�wV݁ �F�����Anq+B)9�>Yp��P�3��So�7W��?B§��y>	�>�h{3���	��3W:�Fá?y"Į��M�d���T�Q��d6�u�~p�KfHD���4��M��6as}��]����E�Œ�$O�]	;a��qW@I�^/ �9hB�mK�c2I���W<T8:Mc?��I|��z�A���)�ȓ2t�&�=A�Ǘj�\�HE�2Q�����-
y�/c���$����k��
�'n���Z�J��d�V���Z�iA��*>Sb���/1|NA�tu��hL`�=��8�V<�tb#7]�gf� �Uƚl�b�.�$�­#%�V�~`�����80�
|jj]/�O�Ru���	��	l�]p"�neV�h|8=I���޴���	��&Z83d�w^�際�R��V1�S��X���e�3t��^��8U3��$���3�ROyr%�lg��� ���^/QY���p��Hv�����fIݚ([]�\���6FP�XL)����s$�/<�6v�}y�w�=�Q�?��,�I	\�&�iq�o��d����+���1>��k�����Xz�dJ��~e"�kV%�̝���4��BT�|fӉ�����W��y��h�D�q���ld90�J�8nJ��Bb���|A�G��-=�������-Zu>Ō���y�QiΓ�ѣ�0ˊ(s��-��0d�������Ü<��kf`3��1��겲+Vf���Q�1[?;À�mrpY�ϕ̛0Ù7�h�:	.����R���HXԯ ��	\���l�1���Y�q9�K���"i��֙2S<����5���-�dC�'��I�-3m�*(�5t4��FGa~[�(��ʖ�c.�nwh�Cg�^��,�A+�� 9"�?�L�"es��џ�����- �.��H �'-}���nhT� �m��J��Q3�鄍���P%���"CO��Y�5	?oC�Tb9ӂ�i��C�8wP%�f��0'Z���ꟿ6�5?��/�5�5�ǝ��-����4[%�փ���b#W�s��[��X?v-m� �
�a�~8�؇Yv$�oD���f���O5��[<?W�&��/�a�ɐ;p�u���``��Z��p+P���ػ�@�d��Ʌ��D��И����j�\~��Rl��d#)���P�M�dn�=R�:�Ս7D��)%3���'b?�k�\��qP�`�������E���{���-�W�p2�]nkT-�T*z�	ӡ�7B��wY�j.F�����c^b�'Pְ$����1�U� )F����`޲I�B�]���H�T�[A�w��X�̌�ox^6���~���.��B�h�ca��XS�[v*������m��Y���ĩy��{Xl�BD�{�<��0�m�Oּ�;.��mSM�-Wj`��q��^�z�=�A�K���e;���5���S��KŶ�i/|��t�`'����5����O3����'��Q� ��ad:{�Ps����&��$v�w^ϰ_H\c��^\g%�9|bd�rm�sB#��\��
H"�	|��0�ܗ͏���r=��J�'�a�Yi��z�t��� d�s���׊E�*��^��(�ͅ���g$m���)�m��ã����|Z!L#�Xy�&*�d��ť��MF�EVd�0��L���"{g�|�E��yb���'�.�,5�p��#l_�>���On���.��>�����'��m��u��#�j��~��J�Q=D�c�2%]@Y�i	�%�A1�)6i�G�;��;�5 ��t��Zg����w�ѳ��]���F�Dֈ�]mϰ�,y�ƌc�vߤ�.�~�l�����ǃ�'���s/X������Y7�<�Ф+A�ԩ�a��3�b�AaOSFK�_ϵɰ�{hU(ӿ�M�����bCT��\-�d�Kb܇�c?U�V�f�b�3Y �����:��J~�R�r_�&��gs�vM�*����5q��!4|e{�u�S��ǩ�j�x�>h���$�\p�mՎTG���>v\�.��n�;��u
�"
N��(���)�6S0�_�P�3�!ӷ�ζ���@���+�5��\hjQ�ZtN����9�g�r�Z��Z��)qD�O��L��L�&�%_����
Y��2������{<�v8��̈́7��)���mE*���#�@�vS�)��ۜX��=���bA����@��8��A42$��_����O,&�Of�Iw�������\�>RJ�Ї̴�}����IE��/�<��}T� �F��vKD���9��=U5�ݒ��ט�g[s�7�	y$=lL��5C������݆���v�?�}Uf��a"]^�+f��)�Xۈ��+�.YzS�X�gɛ��3����ˡ�9�'݉k�YӎWP�G��v�S�H%]Q����M�M��A�s�A�@����1�@���E��ɩ'Eb�������_�uc�p��m��2Mwڧ��CE��#q[��^����:9��������Zμ��{�cHy@�n��]��F?�"y�0�Dg���-ll#ܗ����Y*���#�+�xQٚ��;���q�����o]�����QOl�j����+�]H|s�i���{�y��Y�&A\���n�˕�J)���,"	�&ё(t3���;o?��e]ɺQku����)�.CR>���9�q0~���^M2e�0�8
� `�h�fiD�I�U�y�'fl�E �fϧ �L8U,������t#Ԭȹ3}�ev�?$2�*��=�p@vw�G�i���JCLO�Ӝ�����`j����r����F�CA����'���[r�1C/�Ϙ{��y��v������`谽*�����,�rN%��ҿ#7J�pG�e�z�ր˾�?|w�� �����,���jSJ����B��c ��$���iļ.w�������˴4��J] !Ѥ�K���G���X&���.�J��Ł�Q�2��R�!.3�fx��%���w�m:g�|���P���IX`p۽����,dzp�wqJ9��Lfg�d'�%��?��^"�]��(�;6�s��[Z
+c$-��a��P)�V�+��G;`�w'C�لXBs��&s�n3�d�EZ�Z]�a��5�$^L�{HR�l��r]�
�_<��
l��긴���1"$�n �_?���	W�;�E��'Ds���}�9���XVOt)uc����E*_�X��Zd��L��zO���N�4��'�aZ�x���LH�0�3�3���d	��>���PT�3q�#yYawk�W4S���"��
D�i�853R��n.��{5��~Ң~��l`��#�2��lp�6��8��*�P�9U���U-a���W/JTK=�gH�QڼwW��֒Ǭ�?J�� �� H�rQ��eX�cW!�I������C�o�A/���\�λNN��ӯ]_��|�����cgA%���T�ѳ�Ze��Uh>ebO����n@��������J��3�� Τ$�a�
S|���F#���u���6�ͺ)YG+��MvԦ��f,��l��D�ܻ��!8��TUpx�L㑾k�;N��%�3t�><(~�[0�$�����T��o��8;�M;N�ľ�Æ�����@�+7�Θs�&��ٙS��I�oӜ�ޛ��a*��h�x|�B�䂮Nb6�Հ�4�@�b���p̊�,�DJjm9��R���:{�T��<�x���j��r�@�'S�0�#yͿ�d�E���`�wX�������H�G{��ņUXN��j��ך# �6��|釫pO�
�0�ڟ{8�����m�pDt�E%�de��f�-V��q;���kGup�J���[z�������Iv%�TpB�9O�����?Gm�=���G���黶Z����o[�U�<pS����̤�}i���Jg
�,�K�{oF]��}ȓ9{.��Z&w�'2�nW���@��<�PNS���D�oWM���,�/�K�X)
WI�'X֞��Y'!·9̈�E��Pf)ZO��xaE�I����9;~���k"/#��/��`��d��H��YǺ ��]�
�k0�ik���]�`=D�u0�.1��j(�&�S��]Z�G�)a��N�$)6����\3<�ר�tݵ�xC9�B6-f�S[����NI�'�p��%�c`F��k-w�Є��ٴ25U�S���7d-����k�1��[#����6�r�nl���/)��V(g�8�N�~{h ��ۮ�<|-�(�j�������(g��ݤQ�c\��x=��,�ԏ�5čiս�MD���xz�,�U�68sm�{�r�}�`�l{P�x���܆-�xΦ L�Y�&��۳JY�#�� �1�e�4	Q�NJ~��(�t�8`��:��y��=��5�x��n�k��$������'��[�բ�$0��y��d.>�$���:��ըF�X�^��4H�B�'����$��:��@脰!쀯�i�`D#e�4�Zx��"w���
Bj�y�c�ݖȐm
���8Z���������f����-#ƙ�0�163�t�b��z8E���:�ߐ¡��-��t䁛����[��Q��A�5)`=���v+'X�����5��X�MRz��R��A��p<���(8q�ÔUp�=��� ���ODM�g��,8�f^J��u�r+2G�ȧ�g�̣��������C���U�����)��'�}�kɻ����U�ϗ�4��E�϶�VG5�m�kz����ԉ�l��z�U��7��2#��Y���X��l��Q2��db���l%�͕�5�9!m$�65����!O}��k�qV���H���^�����y#�sN�5��Sy�."�P��b��U����r���*}��ϟ�?+A~B�T��h��Ye��b_+i=~,9]�;w�c*j���&��Ш�.�v��~�M�*��~��i��ߧE˭C�Mi\ICz$��1j;���*3����8t�����9�O���;�407N�!�~�5��4�f(���e|�6���9��G6��!�Ȗ2!Z����}��-�NQ�����'
q�%����������;���48oz�;�*�奈dM��R�Gt�'O0i�/��p�����k���Ö�N��q��ތ'�Η�X33��e���˅����l�ذX����R�"Ą�����q��X�t�b$�g�)h�!�J5E�DN�.���%K^bf?0��&tޔw8Ʒ}>OR�W�b�ɗNJ{12q�L�>�.�	��"�8@�� �}�]	���t(���S��⫋5�<�'8� ��a�{i�6����k��` =A��;�o���pS�����۶;Y��ߌK����Gl��k������/5���85��^��`�ROtGۖ�٦b �\41�c��eg���c��5|��r���G��a�5�� +���f�>�����L��G��:�Ia"��2�������VLv�z��'�M4��	�:�~������8a���1�^�B�U��e�@�#?y���� Q�+nf
���x�d@ߕi��,�k^���P�1�|�]j�����njXy�*��/�,�;D�Ɲ\4�Z��|~�5+5�v��8�Q�r�Q1��TPg_�*��{�-��HO��גw!��Q>��;��~Qd�I(��Z������ql�:�Ғ� B�zMa-ztHf�!v�=9Ji�<�X���4Ť�>Aj.�����A��EpR�G796�nUO�^��~v�A���2�HULRL���<�� ��y��\&�o��('Z[�O*nIɆ�����<4���!F�~p��&?�$��
<�َ���;�#�Z�.���	M���h���FJ���(*�08mg��=�z/��n�d$�Օ�y��?�3��48R�c�zp.�i9�W�պsV��@�u �d�V?�ni�+��N;o(
���� Dڳw,�ӢI�5]��`7�5�*7\a�90evoQ��1oY�n|��l�P��R�a�=e�4U%M�2g̣�%?ȉ
?*�L�c��B��ɭ�C�eAnR��Ŕ-[ ��* .��?TK]�޲��5<١��ҁ�Q �b�c���U6<���%̰�Z��y3��x9�\�O�Ȯ�:��˷:���~ޚ$}Ih_��J]��c:��4����0]C�T�I�G�&sb�h*Oq�'�Eg�Zyo��	�5�N��F�ꎅ�Ђ �)��a�jsr(�uu}4%ufSN�͊�Ӻl:*E�hyz\�]���y�����\n��d��P�j�H���̑03�ڻ���X�2�4=�wA6��(��Q ��3^��tm���;>�M�R����_�Q� %��
Vg�T�C�f�2Hͨ�o�i"g�v<!b�e����¦�X*�KHB���S^p�1�R=�c}أr ������/�A�H1^����4Ҙl�/vg�~[i-3��	<���ʺ�鱣&<ES�S�u,N�[��-�����j�����ЍGf�w)K0w��rS�n���,��"�C6�}ڪ=~_�N���C-��2�Ƈ�,C�&�I���]���k�zI�w5�6V^>pt��Zk���4����	�S�w��|2����'7�^�0�sc�i�iC��N��PX��V�L����P�#?f��!�zl�Fa�J1vWۨ<ܪ����edNX���"gz=NC�U�q�^B��5��Y�uo4c���c6��EJ�u�*���':��Y����_�����C�4ɍ��6_�T��� 磙X)z{��P$�<JA6�:V	&�itc~ lf/�q] b$vɬ.���?�0��dEۚ�#�'%����O�,؆��E���t!ފd��*ԫ0ww�i�Ol9���g(���42�Ũ؄
��N�`N��o
�H�fh������z�Z��>��q 
`���~_r���=`^�B��rg��q��hӼ������ �B
�S}\I���M��򘙠Nu��0�%@B�����������02�,�*pS�so��A��e�Mky�aa�ܿ�.W�J�QO���xΞ�zM��4%�IRŗ�i�Is��:J��5�1�d�L���;�P����ƥ|r�.�pWݕw�1����Nt`�u<ʯ�?�и_Z�!� ��R�
;t(I��ax�-���[��F8�%P��5���)w'7�@:3p� (�\��:�U�d@�f���7iW3�+����@ �W%]r��/~)u�70*}���\��c$����e�*��l5Ԑ���.)�"s�oߛ�����%eBpu,��Q��y�[�d�ݯ�G����~Y��ɳ���+�q�S�6����j�mLH�Y!R��Z��
>�1 ��k���R���R�޹�_QO��Qe�Y��ŗ�*Ј�=�郇P�RT:�uh�U��z��*��w�"r���+�/M��A�J ��>�+c�
{p�����$`˔g�F>]R����wS�����#��Z�4�2ڦ��&{Ϛ���1���-�u�?;m��K�/
X?w��竣�5��G��q}�q���BG�Q���۹i���d:���@t��G	pAYg�:E��)����k����!"�|"z���a����+;�l�*B�M����%>�I������p���e`�g�9\=`��K�L�Q���gtA�/2"�� ���&��i��[��Φp�qq���0��u��'��o֒`�L���{�M*�X@$������]�+	�JƳ"��G\�+!�ތBoB�Qrr�7�w��D�	DI�5l������)��+X.S��8�@��H�k����1�i�p+koIL(��g��R��P>��P�ȅ�ՠ��҆���塻�35N<2g���(�Ϲ����\S�xr���fO�L�GV�TPϼ�_�:)%��y���ő;�؁/N�~f�>�g�`��%R�8�(��me����%(w�_���R�N޴;�����a1����]xȣ�������0l�'�?��ɸ��)�����e]�4h����!�X�lpIH[M_'~�PGyB�7�IC�\�{��n��"Խ*EW����/Xvy����B�M7���$���W����Tup��>��#�1�R�-0���%���]�7ިM ���Ð%ܹ�Kw9S��>�r��~�/����g�h���,��Ҵjσ��t
�6ɂ}����B�[����Y���F�`��b�(F1= �`t�	U� ��S��^{Z�u�"&l�h���cæ�� ��w���?i1E#F%��e��7�l���"*/:��3�A@6��'9����\����6g���s$�d@�Y@������k��c���ɈmI��k���{�;<]�6�V/��Q>�C����4Z+ŅG��O6N�%�vL}����mdm����8�!��t�U� ��(��Y5l�����uQb����$�%n�x�β!v��	�2y�aᩪ��AM�`j�R�u��AwW�C��?��I��i���-0���'/�E�<k�\+����
NjPZd����}g{��Z��,�*�����f��cR��Oe�io�I�{��s���X��%��#m�!�e#^z��>��������)#���i1!	������Ӭ�h��H�>F"�7�q0���ʹ���e�T[v6�\��#j�m���ι��������yb���I^"�&̦1�mlI���+��Ɲ�d��	�����<��1r��X��h?��S����"��v��j��%�9��J��&�����.�yhi؀/I�n�:P#:����	>�Mw�i�/��5)mf%y$s^��	�|wȤʅ�4Mm�࡙��1� ��{<�2�U��˖1G<��@�9�O�v#}f�b$z�m>"��"Q1Kp����P�y�J�}�Q��i�@Z@������d- ��y*ȁ���1�V�̰��l<�CN��%\q�^D4^6���7
d�=xǶ���ȯ$E���qCqV@�U�
Cei�8B�-���6�ז��Եn$��Up����E�jJ�]��5, T��ɬm��n�[�ϛB�zA��R��lL��H-����w�x�ܐQ��C�CFP���pt��I@G�Y��+	�!�ou�;�{c3S���2�߹��mp��L.P�)��NΦ��tz=��ߺ��x�N�� ��^��m��\;�Jחfq}��7Mj̙x���J Vk.���Q[~��oo�������n��kr��z;�H�3F���۵_�iƶ� r��`�{��Ϗ�z�4�eb�֙'��Q���A��io�D�n���K�\w�B�Ue۫����/��qw�N/�$<���)d1:L3��w���9
./S�qu�oBs��w���A=W#ce�6<WY��!x%^/Q�0�
>�	�˚���Dp�L<.�W�T����IM��k���!!�ѷ.�-'٘|��õl,�l�*�2�l�9SN����=#{e�o���!kh\��tG�����Yjϯ����	���K_��;"��N�|�84�B6��jXڹK�n�p2��Q�C����ĵ�?4v�J��?���ĕ���A/��!��"����oY����*���~�����7 ���+j�u'���V[���t�gAVL��=�|�;�=��h2���l�t�Q�#\)~ϼV�Wg#2�����R�\n��ʰ"�~�~�~���a[l���x����ӳ�3�i���W;gr|�W��o};�̿�1�P���|M��IhM��.6����+ʹd��������S;؋4��9¦L@I�tR4�����%PMmeCtCm��{���H�c�������ʇ����p?��3���_m���lt�������Ce����7�p)��-�TBc�I�M�B�X$�3[c����cwS4#sT����Ah2V6tY�"�%[����8q������8��2��P�i<�x)����y�?I1��N�
yA�T�[d�DE�`t������T�����p�����̴q�%_F���U��Z+���}�4b�sRW��.�X]O}�ؼΟ�z<������n�����
����w��L��e�*�[�m�dDnȖN��պ��9�@�b3a|^�0�w)��X�5����#�t�FEYk�����Q$���g�I��A�@U�e�`��s}�*��R<Sy���|%����B�ZS��x�R��v%��w�S����hQA%E^�U��k�*Yc��'�>��$YiU��G.�?�7��\m�i�����T�f���:��DGcv����`�0j$�����������%(q��z�w�6��C�'`(��7�n��z���b�-�J�6顮zX7�K����|��E���B�T?��P�l+J�{�k�W�tg�-�3,l�)���!U�F�o�M�_�s��%-��R���k|��ղ��J�EX���Nݷ�Cb���a��yf��D�u5����H�S�s�eB3Z&�ś8���k�i��L?���p�?},Xl��ۄN��Ћ?o�g������إ���jS{���}f_u��V�,��^�\�٤����8)���1)��~1�~w>J�Q�N<�����S�c��R�����&�vT�����8�uЯ�`���me�ԫ;�F���u�r�ޒk!߳|���媶2_�m�1y�)~Oc�;�"H� o4�}���V�7DP�;0k���-��c -�eC.j�)�H+��ɞY�Y�9}t=>*V��|:�n�fi3���b��u�j��h��@Ž�{�3˲����ڈ��8�'�R G�8�g[�+���ZR:D�0aM��O&h��ݟ�|�4�7�?�:��8���U�Ɯ�����%��t^�a�E|�bR����x_/BSm��:�� 6���㲿���c������|��x]y�ޘ6�BI���~U��S�F6���W���Bl�!�x���ck�̖��56�$�Ѩ(� ~{A���a���nw ��!듶��>e�K��^�w���o/�[�)�*N[긜�ddٻ#ڮͤl�Q���.H��o��\9�=��<��V_�وw�Y��h�Q���G��>zZt��uwt22��m\�i�J��C������7��z���¼/��~�hJQs�����6��ݺ�	2�l&y���Q��2J�w������A��߸,���JKð���\�7PB����R�m6��nw󒠅�L6+���"���~�������-|� �wJ�	��vYq��YԷ��'�@�S��q���z�T:��ik�V��-wM������/��`����g͔����vNfR��Y�?a�y�?�s8��cG��	�E\�<*F�H����ڪ v��[m�j���/�_*�ȝV��y�K2���	g�ȑ0�ܗ�X��!�}�G�X���!&ǐ��<�ŏ�%�w�T#X�_f����T!�l���^?$�+-��:XfOy��l�2����O��@2$����0��P8�7�d��ʦ�ϋ\����8U��A�W���q�诹��*�ﾔ	|	w�A����T[��=q��,946�"�'��c���Ų���
nU {M1
DJ��p:�Z�2=���h��0��u�}>Mu���ꒅ�9��3�P���Byf���J7"�k���c�;��>��G�K�Q�J��C��q�3U�ǇT�C�,X�G+�C�(����F�>\� gR�VRֽQ���v7��خ[~P�ղ�m�l����x2-����8�Y�:X������3T�t��dD�0�\�٢���jx�B�}(o�zS�$Б�]�i&ȕ<B6��`�&�U53��>����I��Ə����p���	�8��o}��4�d�.�|�����{
Kk�5�p��&u�bn�<���x^�X�nG���YAh�'�� H�d�ّ���Á�A�/���.+�u7]�,��B�C��j��c��ǴM_�����s����$���X���^^���'�%S�v�ymQ�(0�@jW	�3ZP���ʕ���6PA�\��g�S]S��^,e�C���F(�V�Y	�9�δ��X#(��Z�p���!�t[��R4�U��?��jmK[_R�:��5�7���2��)��k�,�.�}���SB�?�Ei��� ��0����<(P�ю��eݐ�Ȑ �㽈O:k�f^VJQ�NT.u������������� M�b{%�蝄��ͅB��Q�@O�ud:�Vh�<F_��.��acF��i�?f�FYŇsT*9 4Nmxc�@���A+�u�.w�-�˕?��n۝?X�����u�I�����T��򲗕�$��G��]Q����!\���G�sB�7Y��`�=U��Q88�4F����[7[����"r�͆����{~��=8*/�|��,h����*M��ʮ����u��د0�g\xɿg�3ߙ�xΓn��Hט�? ��#6̊��6�7��Bͱ-�i��z�����^��s�s��FDN���T,m�B밵�>�m�x���8�`�N�C��+�?�����zȎH�%���q�W�x�/�%`���g-�\�אqK�ʼ��"����5,��j�j��@������ш�m2�����x7SI۔�l�T�c�7�����!>*J�OCɿ�݆��G��(7o�'�(�{�F��U��J��ad'ZUNY_R�A�5�xW�7�(i����^�~��&�|9n�݊�b�̰�H�M]��&��[�@O$(�Ϩ�X�ݦ�������L�e�M��W��a���F.e����ʽ�a�<Z@�|���R^�E��}܍����^�_B.��s�^݋���7�2W2�q)�c�S�ʠQ��A�i`��<.��ʛT��k�y�L�75�l?+�g�]�愨��|!7�A�1�Q�̗������6���#��h�ŦcC��$��ƣg5ҲE�
�5�0��.�a�:�G�'��\�[H���� N��ɋ�� ��O���x��%Q���:{PqC�j앍6!-�k���8E�́�!M�Ma���4���y���'Y�:�2�"�kI64�G���+�G;�L�/ל�qC�C'D��.�]���0��1�0�H^�v[}�j{Ae�D
v��r�C ��47�����q���%�,�Tk�`���]fd�?�xO�F0i���i�8:g�J8��2�~i� k�5���t�L����2?3,.�/1w�溨Q�Ĉ�Q�Qhn>��� 5t�@���䙧$��L�b+��h�2R��,�R �	���}`S�4q����&�H���_h����S�߆̋���똠s��u��-Y�6o�6wV�����Ԡ����b42t�m����)���X�D�Pum��#��E���7ox�}��Fk��W%S���n|yd`6�a���������3X9[R���o���g����{��x#����Aj2@*��#R�h}�VB�\u+������'��V�,�dV�.z�Ct����zw�گ&�Nt��^v#����ih�\{���c��� m ^W����%`B��9�p�i�#����$$ @���B���n�uR*����6��Ĩ,Xٙ��DMᯡT5]����}$��^/	x�S�an'�b)"��b�/�m�;
�}�l�,� �u�^n�o	�xH⤒wj���n+ͻ��Q��f�����W%Y��t�?~���=~k��O��"H��
.A�n;�S:H�P��RNE�0�W?����)u!%��{��L���,��o��*^Dg9��[��
b"f9����H ��˾惾3�a�@��i�|_ѩ�y|�e�ti�t����Y�cc j�"��M+��ڮ:����|)�s {_r�~ƵN��s�J��1�>{`��_$a���1�d�g��(����a⸀�@�ٺ	��©�[���H�0�y�n�~�\��{+�����qM�%�b
}o����^ÿ��{�g��zU\l�(���B@x�b`2l:c�-�f0�#pωp��	���p�9�H���B%�$���{���]��#���\����q��7I�b$HD�� �i�d&�}�!�)��Kr�r�&yaŶ��
3�j�}ef^�:�v`Èt۪SJ�:�\�\.FX6f�Ze.�	�ͤ��v�c���g��P|�V��`�J{|5����ӗ'jψ�<�
�:h��@@ �o����挰,����"`^bG���/2�h��P����>51� ��vN�{aOH�O��6�`e_���ܓ#�18�(`��M��"u���%��eEzɄ��%}�̲q*ZUJTVŶ@$=\�j��h NtC����q����eOmRSj0���A��ݮݠ	6��1vS_!�Ci#�vU��ml`��濲3d�b(��k�"\pI�ͭ��8�x�v}θ�؊�������8:s��+/��5�Ѵ�-��6��4�iy�5S�T��!9�A�zx�Q�2��m��a���[Q�5Ɲ���|���Xt	�	F���_̈́�GI�xL_'����B�T�2�c��6¨G����C+n�?�����۬L�'H���A'�o4+;4���G�N�����1�R���U��Y�ϋ�Hov�	-G�<U�W����J9���~1q0$l	�9���$�Jn~����!���rc��Iy1����?���Yӧ�6�;�����s�r�^����tٍ��-��;Ňҩq�3'���ΚM��}1a,��ϖ<N��I�*d��lH�_8���iH�1��n��Y�Y?&�b��m�5��Y����,�'�x>�;B>��A�킮,]c�Q8�_��p.M���Qi��V�$�j���6HE|�������8�������?�`<��|eo~�3��{WA_�������`D_��u��b�	�����{#��_�q>f�%�eK�4�^N'����ۃs�bb�7�J��_��M����ې���m7Fn�}@g(�^r�Fi	���$�|��i�bK���[��t�'A��I�(����x{-pv���G_���Z�����������T�	g㿦D�C��%��c�7�	T��x�>��_tr��%p�~���1@�\�n"/�Ε�j���#��6+-���U[R���Z�W2K5�uq?�����!j ���ewX��5Uwbd��.\
���TȡXc2�	?l\H��5�I�$�}f�J�KD^�TS.����d�(�����.����T���L�da@��3�1H�`R<F�;z������m�|^�7D�B'υh�D0v*=e�39���B�T��J�`$�͒���$�G�+$���}�q%*_��T�5u5��͛�Qdb����f}*�� �T�NZ���d*�:�m(�5ǲ$G_�����m�eK�p��/�hH.�x����s��w�=,,����|j��i[묛��e��C���@-�A�]���,ڂu�����t<�(�Ww��.�i��x�T�������m09�/3����=�pX�6�&̈�O�����/_�8����ꘘ���<��e���r����
Qr�{d1+q*�7�=����і�G�*�����@�j���np�v�m�D��c�����5�	 }��8\^6�2�%j"$��ΐ��#m���]� ���s��Il��1��h��>^e��('��ԜWJ���u�0f&d��1^���5�Fva���[O�H�d�S��ɻ�%�w�<����Q�R.����(73�z	����n��;0,Ms�T�^��'M�98z=փ3�b4aqp�-ȉ/��7�䰌sN)�u�����B~HFl�vJ~�
cs�u�41�``�`�T<����#6�4<���0)+��F��#(�Ҽۊ>�E�K���:�I���W��!�?U\��ἎY����s:v��K]�y.��D� ����s�E�~��7���~�W7M.J5v���j5�Ri$Le'ɴn7�b��m�[��9l�1�4�a�c�oT��oV�Nq-o�e�(����S��&�bc[�v1DSik�O����%�2�M?A���'!��rj3s�{Z��,���fuA�Vs��b3��0rЈy�r	} ��[r�&�~q��n�^D�+2 ���(�z%:�˴���e�@*\�n��)S�\���W�w\f?�LW�����xΧY(�tnLY��^7Y%�%���K��Zm~Ռ+����c� d�]�Cn���I�!���@���
 �Y/�@�ԁ���:3a���H�9X.�7�J�����_�Z��5 ���d�JP��d�����#V��Nf|�%;���僑|b�&l��^}�?��E`���oT0����J��_��L��r!m�n|Z�p�`r�Oud���Ʌ�;<i$�ѦBл����{E2��������[����_�����I�
�n����Zw1���32�Tѿ�ɷ���ԪO?