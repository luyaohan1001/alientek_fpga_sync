��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G�['��7Ⱥ��P5K����v�k��8����H�V@[��;Z����bX��Q����jF���TN��L��l��:#��+jZg߽Ԗ������MSY����!����<͛?�M�ﻼ dc/��al��4��`�ؒ����i��e�{H)��	
V�����O�h	�S]��1ֿxٔ��cB��}�9k���R3����M#5m�J����5�������ىM��Ng���G�<����Z�"�����\�U�]�a<f�)G\����5��qG4	�C�vJ�&��{	��5 -m,�8�kK�p.��,V�xy1!���4���[je*{��#��7���p~T����<j��7��v�;4u��'�?��^`�%4�P���||d�l�f�+��<�J��'���fO��)��_��cĎ�\R�9�m�������!��i�X�^N{Nh����U�p|�Q$���^?�>kF�."b���d���3O򕳜B���uq ��r���ǁ��x�f�T�0�劉ފM)R���Ր��	�EEw�8������d/��a�<3�ԑxk��J��W5� �-r����~�TMr~���q_u���ɬ�I<}�g����2D��X��#��I��VЃP�?-�fun��������C�_t�� ]������,��e���f��v��i����6'�8N�>�')7�
5�F*5of���#/e�40�znx�d�ۥ�~��
�f�AیW<��,S#�i�)�᠆�� �A���at�wA̍ޗPs�*q������`3ɤ5���Bu��K L������3�#GGӈ��	�<�Z9}"+���X��2oL���6�SKtOK����ӀͻL"Z^ݢ�?�G1�V֮��E|c7�$�6<�4��3q�GtÝ���k�?�&��[�ZhC
�&�s�������	? o�FDiS�hj���g@+������4��^�A0V��MX}�?�veT�-�K����c�V�g����	�7�� ZY�t����I�C�P6�c}��'�a�R��x��J>��u�z��Z��8��/]T\	���W[!������κ�:��0��ˡ��ν}+��C9��xCL�L�������H|�҅��	݄\�D�aawd0�D,�Ða��_���(3�Vb�'�����p����N ȏ���fȹ���_��yi^�!�(]$�jdcP�=��b-$�2�}�bQ[�mȋ����4��*]�rO�R�GS�38k{�@��sM`jt�]H?�a��w�o�����یEED���d�"�j���5��x�r��]�&���@�jS"r�sS��!k<�?l0���/��W�p��߫���p���H4
Lx{�=�4 �.����?t^�%l����\ш皜T�,!>�E�+���儛J�1����t ��_왅)1��q��S*;!��&|ז�����͈)��J)�>UӜ%��<G�6y��f�
,E)��3�hT;t@�c�#�
��V6HP�4�dVlh�=�T���N�<�+"CMk��U�8�p�D߉���#�t�s��nu��.yc*��BD�{R���iI������vnaB�&�b��0���n$�3�$��)8W��4"y@G7��P%�U��R�C�,1p�	 �Ŋ�tS�e����P7(��|�b�褾�����p|������6%c��߰��^�R�-�+ 9�S�����BxH�IH�o[>�%�u��|Y��N�S\Ҙ�_�&P�*��7h�s��2�����˂�L�~�H�s"���Qΰ�\��њ1/c�/��7�C�h�f���a�X �����÷6�	>���qOP�4�A��$!R���\�ZZ6�ΊՂ��j���B|��ƃ}}��G؂����a�{-a�$$0V��ms�B�9�*T��Ii;��r=�ɿl����j�j�9�w.2�_���1�kW���f$.�.wu�?�I �dD��b�j4�.���J�W�ȑF��KMF��OӶ���'VYH�
�'�o����	�L��d��!�����k"����1�,n��#d6�Ħ�{����;�s�\���J��S�m����Qz0�s�r��S��@��jug�p�� ��Q�7�ݼ˸���DMob�u��1{��4�
�?�� �:}�E��r֒�}tL���:L�����i����j���Va��YO{fE)����M9W�������S��h��ԡ����6�So�`�D�E,�
�����B���k�#褓B_�Tjr�n:L�wYG_�W��]��n{��2kyU� �@	�W��u��v*U��P���#�nCH��q��B��9�w]���ʛ&Fq-ٱ�󘸻��5-�AʻSX�t:��N)��P�rX&��^��1�3~��	,F$Ԫ �+Kg�mp��6�N��j�d,�­z�_���	(�k�+�Fc7�D�I�M�5��j�W�槀c#`0�l���a�h��䒳_:�2Y.��	�����FSKTͺ����^���C��EEj�̹�PO��V��HT�[�S�8�O��>����>��G�8Ծ� S��{�'6�0����]�ۛ���^%��7�`ge{�6@�c9�`)�����7���n%f��HQKJdx����M���b��ᡇx&��Uh�J�i�]����v�u鋑��t���L�؀m�|�+�խ�߰Q�� &	��_�[�*j+eXcӕh��ٽ�h+�vB�@Z��*7���+I��r��yj�#�f��^��aX�x��Z�0&(6
�4�/���~N�P'�% `9�}[�K��ԗ��0�w_ۮ��	<?��.����ϠQT��B�&��g�	��iq������U�K�,p�΄�C(��V�m�آ��ƌ�DQT�s}�\[Z&��Gor4���_�_�j�%�P<R��AI��P慧Ϟ@�����!���ʲTt#$	��:���O�x>������������6؂�!�.ԫ����`�?C��v��*6���s;�eg%Z*$'���;o߈�sӦB�?hDb��S����ߤ��8KY�^ϸ8��16�yђ0���b2�>�����s�v���܌�2��`6QI��:��X�>RUv�\�{�ٝi�+q13�EBG�����"�L���,��o��K	qw�f�%��H���g$��?$aދf�|_� �����X�=v�����dd�0�R~�]6�{���%�n��B���f�}9!uAxHI/��${<Z��G�ļhlE��Vy~nʴ���1j)�A�P�^�'�SP��{�(
�����tZ���_^�{��sܦh����9o^�9"��e�TS]*-�F�!��-���(���3���Lc⚺L��ԑo�C��aݧ�4��0����F!V����:Ca$'bZ
q��2�."%.��z턴���������T�ψIx�WT
�A��"*��D���w�G�KW>t�������t��� LRWv���՟�m�MN�L%�"��_y������$�#�8��فB-ejP�&Vw�"Ƭ���KI��|�T����dW��R*Af�>�\%�@��n-ᇤ��^�.����T0Էc?��u5E$�I���N0�eՄ�Q��Q��."���=�tb�h�y� ���	�]��9���_������4��oU����a>�E�LI&=V��ɠ�a��Gk�����l	H� �C�ܮ�藒�Kh�αOb\�^)+ٴ�elɂ�5k�F`��Z���0��)���h1+���Ѓ�tQ{z��T�BC��J�1d\�LJ�>U�=پ�o�E4>	��`I`n���c[��>�7��G�������W�!]�u�oh�c�C����	�u~�^�S`"����X�7c�fX*�u:�`ð��s�=����K�F�� ��>��W�c�P��bp��o�ѕ�?��I#��qj���c�ۍ���M���v�@{s�PI<;j��*�s��ɞA�N%�m7�D���%H=��4�tV�:�}GCASi`�6/Ϩ(�N��ہ�~wWN������M�zy����T��R�ɧ6-�n0�$:`��mm:��F�����	�?�D�P_�hn�E�R)�c���p��ɏ��-�ηz2��,&����_���M�	���y+�-�ϻԙ�/�#[��uh����8�\q
W}ɻ@����h�3Nr����9:`�����'��%�ck�K���!��Y>x=�%ҙ)�5^���q-��NGہ�[�~��C2������&���L�r~�O��_�F�R8�$��gQ7�i־�C� ��Sa��2Ay���p�9��
>H�`vMę38<'�d�Ύ����4N'�ʐ >������?�����De]q�)�/;��Ẩ`�º_�k�V���R~��{��wi��R�(Z���	ӻn���x<;���B$e-e���	I���i��i�c�D~��Ь��*����|�Ĩ�S`Z��搇G��JD�)�M��w�&3	�,.���R˝��4��R��4)2��*�_��{���m�0�����`�9������D��F���׸�WD�[R���_�q
�Q0uڱA�?5�ö=�������	���N !Hz��дJ��}XÐ��P9��7�pFY����<�먹����6�=�(K�c�e�&���c�U�$�����{"X��W���ho�g./�f7��\�Zt�כ�P�-�����m4Rp��/�Sg�����-�Z�1Sdl�߇-󄞱�w{�'2�z���ץ�湙,�z�/e �.PF��^/_�D���.���ʣx���Y��z�����B���������y�R��� K�ƌV7�)8�:���w�6�0q{;���^�R?cҭԿ� 
����qJG(�����u$�rQy�(�` ͰL$2�������J߀�BYH�cj�ð�D�T)��G%�?��
���Q�Z̩+��$O�>EE�]B�CU(���|ځe%��ĦF�Di�C��U�9N\�E�y%�XYy��.(V�����lfr2�����T�1"G���V�:N�H�ڨMMJ���r�@��]<'�YT$RWg�w` P�}!j�Iz��\�<�"p*l}[���h�Ymt�NWx.5��Am@m!�6����ʚׇ�q�c6l�;,OV��#�7C��������u��]��@��Kj�6N�22@~�r>���l���^���[�@���ֈ`�G�hJ?��c�����Q�-q���*R`W��LԕT>�BƾD��!�^J�?�@��l�_�OlS#�U.'dF$k��zXEǬ˭a~xK'+̈z���.i�%�*��i�H;�l9x���y����%�8�G��������9l���V�]��T� ���������)V���-!?w�6ї�^��[��+���;�
��s�(�bׯ"m�s���*YQ�S�Ȃ|�y��(��)���A9��c3��� �{b�d/�e2!�P���|��K�a�qt�Q^��m.��Hj*��nC�?��h6JJK-������Zʔ�r���sy�"�uA�	�D����i�X�ߗ �٦8�_ܿXtu0E�Z�|�`����u6g_z��wI����-�Z��'�S�.c�*l=�`�6K:+a�^.a�p!��:>/*���(qs\|��vw�k2s ~���(�=�mY=	�lthΙ{�y|�4Z��x=��њ쥔u?�	�����<0c�7c:tV�2�L|�e�0��Ĕ�}
����g�.�\�� �?%���!���
±�8�&��Q��iwķ��Z<[�;�ݲ����K�H����i�Ͻo�����2X̼��H�H���r��Me0j�a^�"�-�Fc�Lmʉ��z�@�x
��"N�6QG5?1]�$L�k*i9.ZщXq��0�@nE�2P
��� �Ωݺ�	��;�6\:�a2nqp_!Y����棲���97�����,�"��U��]��  �뮲U��Ty�H�����'��`� d23�@���A'�-�3�	gQ�f��Ds��,�ˁ�B��N����~�˰������Y�����<��*a��AB �ٹ���g��FX��'[f�d��ʘ����������\c��(]M*)�&]w��;g���w,^KC�Rg×�E�n����|f��~��1#��z&}[)�`,Q
�>��#��F�P}�
�6G7dqV����R� ����iC���� ަ�8*��it�S�m����D����`�G�ft��t]%Ȥ&"�w�P��G_��-�pX��9����J��?�c���@j��ﾟ42T���I[@���nm|����Ҷ�0�JUW.��C+�}F=M8,>��>,#< ע·q�>���{�^��>h��t��|۳�Y��٠���eÃ���æEs����1�_j����9n�$�;��L�C5���l�*���F��~��~:��iTK��z5bQ08�'�j��e�YNKA�®Z��œ�4)����uPu��R��fb۫X�Oy��^Q������.�AT�w�J���t�sޙ�\@mB��PqEN^q���͙oǕ׬�[�ɩ��,h�����}��k��g=W�KNQ<���C�n�t]m��ik*L����R�@-Zܲ�8ui�������������O�������e�uD�����8�/lM�g�k_���`�+̆b+K_5��r��9e�o�e��۝�/�W������e�&9p�jkx��b�}H���}c�yj�rj��T�L��Ql�~����<�a1���
ȣ'3���k*�N4�z:�M����OE�D�p��|���3�{+��TY� ��} 9�f����9SԷ�P2�q�R׋��Q��fZ���A?�� �Gɕּn3\Q�����eu`�G��޸UUT�fqM?�7F-��U�3��IC�����|�r �w�|=:��7&G(NeT�ko��aO�pƼG~���9�W@?a�!"�{x9�c��T���N���t���s�ؑ��)T	��HKH��m�������q ����,��~��=��7��`�\�~y�S�2�Z��
�npĥ��p%�<x�-�FJY*#�/���tk،|jj.��4ˑ�An�;�fy�:#�[ 5�m�5��g~���WZ��3#J'�G:s��k9'0�� ��G�C��sD�R��r<Dn$�C�.�IӶv�;K�M��I y��p�`����Ya$v#2<e����
Sꆴ��6,�i2���
/� ����2zF�
|A�m��hzĖ���W�$ �'t���zOI��%%���	�F�4Vx��5�Q�(���z+��u����j�e���˹A��L�	z���'��V��h��v���g�"�ε�z��SPhM�̆���һfß����\N��|)�NE7�-��)���!@V[}��{o]���4oȵ�1�x��p�`��2g�@�b���,��1s�8��T(��te��Zq�gF�vz�r_�=M����c	#u���ym&�1�.�[ ϱZ���̷�OUN�#:��TϠK�P�o���,J́��թ����)%yp�+-dX�C?B1Dm�Eb�����ct�Խ��@�S���u�0<���zy=W�AaI���ۆ�W	��6�3�5�x�"�XW����N7���b��dQ~a�c��K��7nJ�jO萭W�rƿ�oC�F�Y&>�{҅�k�,�s�6�4Т�f�(;��Q�w��R��׊7��[2�\�\ڇ����&�zs_Ѝ�����m"�4̹i���yI77�K��X����(�r%�eTm���,�e�Ms�ۃo�X�'R辧
o62���)|n�f�7��K���g�����/^M~ơ~M�
	N1�g/W�������i��K���ct�.+�Qo]|^���9��t�5�N�e�@��̳�3K����mo��!����b��/��se�|�r��` w�ZOqt��]۶`�����+���6��f�Ϝ�Y~����=^I��pm��~nlr*| A��%��??���
;M5.2��h���մC�1%n�r5ITo�X[�ؓ����^c��^7��<����2�t�>��#�?��E�ۖx���3����'K=0� ����h����UaV�aX�,�
m&9�D�:����F����L�C�d����l�)=�&�Q�� XE6�j��nŞm(.�U�g#X�a`��*��j�$(����+4C,���P2�Zu��͚oQL��؟_�pyN24c�'�����P\�"�X�3r��==���ؼP<[���x�'r������L��ߛ�X��sZInhB�1��I���\�ū������}A8m�,$$?ēlJ�Jr�k����	eKWV�G5��"�X��������h�5i&��~{�L��%v�BۤR������MMp�����k'��#�_�����}�j)>�v��SGȸ3|h����	�D׫�V:����=CBUp,��z�-���G�d���QV�|a	�=����eM������G�`��C��E�D�s��h�uqE7N�eV�7�l�m�f����v��?϶�=M��re���Or��D^/!Y1	����1���/\�k�F�Ρ��<��'�S�@��5��8�j�����\a�f_Z2�`�^��IȎ���b�|	��I����_����E����.ORȜ�4���0�K<pr@�/w��{��Ї{r�RIO��QT�x�B���9��m��μ���R���g����w.=AXe�����J�6��M�JB��H�AS���.7=�u|w���8��g]U����J�Ɋh9�"� ��S��,Z�,c��sP|\�z��D��?G��7�����˽�30Aؐz�4�1j�ֲ.x%/�nr��j��+�K�&���|-�a��XKM��_�[�T��{ ���)cl�ǹK]�A��R�k�ه����h��G5۪��	��,R�D��|�����"�w��kA;g�_��妪��`h�Rm��ū���R\>$�)�.��P�7}�g|1��1�
{����+s�.�Q�en�� %��j��Ρ���W[�%���)?� ��R��St"0�{~_��e�Ev��ɉ��W�k��S\�?��u�'@�@�ܖ�)�I�߭�Xu��Ň�-��ȝ��:/�,���j�݅��t��}��l�}Ƈ�*��T����9��J�|�J�ܒ?U�9εa�<��H!���'�����R4�RC�L��#���"��(W�r��RB��]�ƅߤ.yb����ԕx�=���
s��3�o��TA�#�TdmLF-��Rm%�G�|2�9F���������ɯ�Ŗ�z�9Hy/�	�#v����Ϗ�ɧ��%� ��p�d�ړ�j�Z˵k�C~�q�=�,9�<u��y�m��P;��݌$�U���6�2�Sy��9V�_s��y青���m�"D������|�q%�Ŭ�}P�1;�w~&�����4�	�Qظ��n��F() ��������u;g�7�V�(٬�o\4����Y����
6�¦�z_C
XP7��IϚ�T��NÖI�-�������J��>!�-|��*!{R֐��*���ZK��%��5��H�I���l-���f2�4���+�i�&'�����Y��I>��pj\�D�-�D5�[�g�T�iut���h�����ug^jD_}��+�|CO�N�S���-F� 1r���Tټ�1�t5��12A�k�����D���mD���R
�/}Bf6�gQe�4�2���'u'�%��a�y��e�=R(o����ƿӜ�?���q�.̳��E��)C~�Y0;��T�q먰րXƢwb��Fp��q���En|u#��d��K�C�`�����zwA/x��o�{RxU��������S�0���I*ȴ��B�rS��\�(K�(P���C�H0��A�kH}��`>��0˷��?мC����Ԟ
C�$*t�@/����<�>�$К��"�?U���j�D98����!l�)v]"X\[��N��޳w��:�'����$�r>L�HcI��@�7�$�L)����P&���j��R\b3@����C&@��#<~:��Vţ���s���Xn;�c�G�i<��<%�]{�?�l8^J��E��WMiuw?I�̏Wd���-dt7��U�>����7�'�K֋2��3E�*4I�:�0 ��#�@ŞK7|��͇�Q�� ō��~B��GT^�.aڹ9$3|�й�GUҒ�B��!��A�h�Hc1/��|v5�������*imF�FWV����m��2]���K�$p�6��l
�ք����w�3�Ⱥns���*Ý��v�~��U�.�4N�頾<Q����t�^1R�y�6ɘ	DX�69Ve�1���<`k�ޮBd��ٞ�RN�ޮ���D�*�s\�1�A?D�"��п
b��uca���7Uc�-`!Z�+��L�-�u�s=��sOK�mZ\���F�\qFs |���{�,<��`��j��Жe��Θ�R���3��胹u�K�$N�<"�\�-Ձ�/C�t�Uiu)�U��z*�{M\���|�q]�(W��h+6Jܲ��C�����g
��������Ub��@����EYP&�:�W0�Q�Tu�ڡ/�V��[a�%ٯ��Cgp+�� ��z�<찡��
}����\�O���Q/)���'hX$J2J&��Zs#�cɊ�,��c���e��FR`��F�	
>��.̿�<o˖��]�6ޯ/U�?(����>^�A��� ��&�Bz�ȩFF���I��~�^M��
��L��y�*S�a�N,����O�ύ�a�^}ܝ�M�,�`���Jd�����tJ+%�̘�I;��Q���ƻX�B�}aU(�m���YCB�E�E��(Ͼjȓڵl�p'�W	��9>@5�j3��1�H8����]�R��
 �G@K2�Zzt{,�3��gT"���!�o�P���a;W���g�3F/��.�@��޺��95�`����mF�i�#D��w��"�qA	��K�W�.2�i3����W��sp��+S������MDs�Y��H���n�*��o�{�Z��f��r�����:����C^�� �$%�<��d�� *��V�!9�\�VP��IB�?IƆ����y��!5`b�f��|�����n��ݞ�Cif�$M{$�Ym��W�l�zB���Iu=X ����RZ�H�
\���Z�<�P�7�&ç�7o8Hk���f���W��N���0�4�Z�dWN:J��D�9+Z��K[�y�qhD-%\0�� ��S�,y��Ytj���z�qz]�5YT��j�)&�ߐ�p
#\+��;�j7�K�Q��H��� g��Ӭ���H�I�����ߵ2h�L�~I���	�1HW=��:���[q������O�#OO�ZA��]Xh���v@�����,��-�+س�#���s�#S߆�
�	H������=�� ES��=y�L-'��.��xQ�w����nĽc�(��	���d7Њԗ"|_(`�������Ep��ȴ���ϵ��
u�Բe1�?yR����|*	��kЩ�e�m���LW,K���զ�8oQ&(�F�dQ�����3�ժ ���'���o]�#�:0~��2䧉�>O�6=I���i��)���oٓTG	�-#656�3C�O�M������W`�U'��W�lЏ~ȁ��T{?}m�N����2��8Sv�i��/ŧ��׶���Uv�����M�.,&Ŧt���0~c;��An�$�e��!Ηŕ$7���~Mm�D����Y�_n�������K���ۣ�lW�C���D��t�ƾ���T9�j[O��4[&�Ն\���Ð��(Y�$b�4�Y)R�/�o͢�XŬ��Ɵ�H՚�V �箲��n�%<bj�d)�vf���X>�EE�3�ё?�%�!	��2�┱Iy�^�m�*�d�.����F	���e�1�àr"�����n�f"��( -}�ʨͶ;�Wi��5l�3oB�i3'�M�;�t1���Պ13��+#�%�9گM����/3�%�������~��W���2v�A��b݇|�%on�����e@����Ӛ�� �0D��a�\�¾�Y���v���u�F�ہ�v��.f�_�3�1jd[!�$�8WX�����V��������&��r}��YJ���Mna���M>5��*΅�-�h>���r��h`KN���Tu�gh�A�Q�����8	w%�`#�K���t9��Ӭa�1^�Dc����UGN��70�ɻ,fHz�ۧ��eo�x$�RT�$w����0\���ݴ���=qP����XV*1�c��5�%��b�vO�,(�P�\�C�X��Y��x�r���/�r��D����Z��׺��5̆������ul�	��vL��0���޷/2[͜nŹ�GhN����P�᷵-�빘�X��m%�����:mn띺jM �.���Q"QmmBL@?T�s[�-���Sgb�U�ҡ�݈]�K���{^��Ʈ���%$%0f�������CX���8�kԦ�״8�F���kP��ڪCa�X#��
G��Q�CA,�U�����}W}���Mo�l�,�(݇���e�E�KE>���������	��cЛ~~��(��j��f:��8�;��S�Ud��,�7������8�K䞡MW1�'���BvF�Ñ�щ+�݊���bL$w��G�d���(�8T�o&x�dJ�P�|]��xx�9~>����]������+���ͮ��8�"�4���� �䟛�Ȅ��3|{���T���a�����P�֠����o�(�v�	�z�~�A���X�+Q�ӳ��1�Œ}�$z�� �q{�R�c]/��i�EY�I�����G&k?��<�z)	\7��G�2�D �s�uf��7HR3*�K����+�[=~��k>��~�K]�kLT��Xud�-9�x�{yQ��y�#e�_;օ�=�r���!T�'u�ɈL�&dP��׭c�
�7�W��*�����,�o�"�����7�$�g�Ck0`�� �&^����頋���C���xG{�E#)�4߯.y2�P����(%s�[�@E�|�ܰ��@�(j���j�������_�)�c�f�@l�9s�뗭0�{�y�;�{�|��>Մ�:��I:sz�@�N��rDE$\��sR�̎�B�dm��N���������������,0���Kmo�.Gp�C-^W�dW�L$.�ْ�_Uq��U
�}��`k7FF;�_�mCN/���c���*�$tx����T-�(�C`U��8�{�{"�.}����܁R��3�(ag�N�^+gv�8hϤ-5��\dQ��O�<�l��RF�mC���g�e.qy�ЦݛJ�D1�d�.�;��231 4I�TM�aO�<S�@8ܔ��
Q�[e�}q�]���������uKLuRo���K��r�nI�܆�������&:�=s����Y�W�4�͚�am��"�Ke�%�����Q� ��!B�H�}��1h��4q�TOҚY"�"���7��q��x���$ȃ��(�4���a�_�&���_\qҦ�l/��#�j�oADb��
ʐ��5�$��;+:�Q����A[�?$��p�cj}���k�R��5e^i��>L���ia���Fi�c緭�b�[%}�s3�v������U\7Μ~UeRr�}&��.Y���L�g�Uu���ul7m9�ti�!5�y.�Z��J�VJ�z�gD���<�ԑ���4�P��S�_-�>�����J�EM���4K/����*�
efbJ�*���IMI����%8�ɀp�P�O E�f�u��W�V�����s��y�S;���3�S���B�K1�O�����A�NUH+B�n��6��ן�Q�yt�Ô���:iA�	6�XiR�G���eMaٝ�Ԡ�q�J)��+�J��$�_�A܆�_Un$.]]mI\	-��Ô=ňu-��������/SmPF��Kn�{�3�|��

<��B�����p��h�aa��gi�&�hAH���
'uY��?��e7��Ya��@By���\��߫��%���<�6Yc��(i�@�� w,Clʟ~����!�n�t%���1��B�>������Z���k�2���p���)�w���ݟ�d0��Yz�qeUU^�5�A�s����z�@�d^��P�I��ݤ6^���j?*�VG!�K�ǽ���;��3���?ѭ��G���o2�I��8/��$�s��c�]�ͤ�p *�u:A��r�&
!3�ۺ��&;�~����5	��,�SJ���E*��G)~���l�]���9
�M���X#�jq �%k���5�=��]�E����hwu5���G1��4#�E��\/�t:1��6�p�-%��Aص�I(�O��-�b�n��c��Ga���p������ߠ/��9�^eR;Mڪ�Y����]��ԿpZ�a� ͈�aȍh��~�,YQ�E>�E����F�k?��G�]����U��{/m�b��:W����A�i4������`�*��߳���q�-�,�?1m"?�E��BD�˾Hs��n��	�R�ޘ�÷M��~lL�����V��1��g�K�-��pge�T?o���Rs�#� �I�F�u<@s�`'Tl�� �S���!c����3x��>��"ւ���p��9��H�B���W��P@������k7�8����(��4u�JLx��X��R��2'�)w�Rn1������]=�cJ��&:��N�)O�k���U/{�^�׼}�g�]vo@l*|w�W���íuSt: ��,B����R�-q�-�g�n���\p
Hy)U_�<F�A�咒|��gx�x��el��.3D��&}�q�!�G~���jc�2�� ��q��0�o���4�%�ܱ��E�}�b�;E� ����#H�	�~����˺���6��]�����th)��j+�(�j�"��CvaTɣZ��^>8}4��69�M
:�1�&L,b����i@��=S.L��5f�t��q�É�[���\q�ٍ۳6���<�Ġ�<�(k�	�&�+�#�W��L�Y}n)�W�Vk�do�|���+W����ɤ�	�!�������C��^�l'S�����(�8�����Z\~�����[O^�QR�#d���� A��������d�Vj��IgWTg��u� 8��D.L :<�[ra�'�^��������e'��R�aI�7wZ�4!\~����)le�aq\v���.KS��qY��ϗɝ��0Z�ExW�DM���<���dVƀF�~(�����о"H�&�4����>n�͵�k��ך'��m�=��9��I���zMց���j�c~k�I3/4+��G��6�#�wV��Ȕ��M���㞾�6�6���À�WSo��"
������h��e�?�.��'�뛼�8�o(T��V=�c,]���F�A���v�Za�51-<� tU2,�W�.��02��E��t���]ȵ*Ӭ+�'se�/B�����:�lg	bVǦ��a�#5��`�W F�̮���n��k0��zo�N���&�������^�G����2��,S¯�8H�6{*�7�(�Z���~t�U�ܘ��T�o�I8�g�A�S4;�	��+At����$�^�
R��P�0�"��uV�۰ct(��<�f�o
�h��|�Q
���!7����T��J�/��T�FTH�!N�{�Ag�����;׷~ ���J�[M��k����w�ˉ�5�_s��ܔ��4o�g��|O�.�� ����-��=���W�|�<-cNVG�24�i,�󳞕)R�����9@�S�a�jg����E��d�ňHfN%Iv8�����KE���VCEI����!?Q�ַ����ru���~��"�* ����� �'K_t��c��O��� �o�O�����X{$�e��_J_��N;|���͠���d�Ѣ�o���q ���m�(���J6lY��{�)��~Z�Fꄹ�TA���Z�Q�B�HZ/:�9�d� �A8�3����hN=*�w�T����7��`�m��$�Ā���U�ɔU�O�r���b-�R}B���1~���NR��$��>����_K���5�T�V��+m8.)(���sq?Hˊ��n��Ykh��/��0����@�2�
Ă~��nI�6�4o q�TJ����-,�I����B���9}1q6��'�Ci/�F���>@z��#M�(hG2��!��Fw����Հ�~�c����0B�K)G�h�5D��*���MΖ
��3~�[j�����C$6r�pB��6A���f�>t�}�Y�)3Fۉ҉���VaS�i�%�+�ӑ*��j���"й��S���H��>�d�T��ҫ�,%� ��|BMdY���NXO�������x��K���5�O0����,�xf �!Oa��@��C������
t�e�jB�=F5s$.�H�՛�46?KVC���#�� R"��}��P������C��J���!�}$}�J�"Х,&�L_P�y�ǋz�.�\;��ë��	����Y���vxӺ5�S�sƙh�_�8.��("��7���Yٽ-�����a�V��
)�$�J�<'R�7�'��^,|�q-%��YO܆H�#�I�a�v2�t��H=<2`��5w���T+"$��R��{�T��|v��-=�����x#�_^Cr��X�����Rh������5ԭ��(�$H����höCX́��ة����H�z�y{��L�bW �W��������p넘����p^4��5�Lv+�*���v��K"��24�ĵq�	�!6�Ŋ���*g/�q������m"B9��/�`v�i���n��'}ʝ8��6/�_l2#�����"�\�p%���d�U*K��v�����6�qp"��w�ҁ��t$�=f�`�n�Y���-C���C�LN�=�W��)]3���>�=`� >7�<�� �
i��ZvZZ\�䗎W�ٵ%s�T�C�5&~��D#	a Tr��m�^���	6�������*�����W����l����U&�����#�wA��Ip^�-��!ל�3��NޠQ�S��9�N1	l�pJ���>�C{�,h��wJ��9��_��0ڞ��,�YF❚h��%�i�q�ղݮy��&U���b��T�������,c��?s��0x��2�5�3��ϣ��q��Ԩ$���^��5\��v�u��6��#�Dm&S�� ,<f _]ѝ����(��w��y%^���eE���=�M�"b��G"�#��a�%�.�`f�p��=�y֖`�_�4�l-�xl�u̇�f��(�J�\"[�,+�Yrs?��{|n�����~���!��I���
<4Ҍ���o����튒"�BPaU���EJ���^Kdf��_ę�!�)P6�aX�L	��/e����7�/���'߳��4��s��c���R٦G��F��]����8V/8��.�1C6��ۀ��,'ܶA���%o@(n��]l��/�ி�����T���Γ�M\��8�e���J�9�;��9D_	c��M��O�C��7��ꤼ�;�^bk�<�H�iK�pJ{4�1�L��L#1gW�|c��?]�cp9�f�/wA+#����������5�K\ت��E��̮D\�.�*N�^n�_�S�
uam�㨌�\%��|5���Â�Se`�U(�CB���Ѕ��ڋ �N��k��^�5�g� ��4�'+�+?C�88�]t}{(��N�˴���7���qE��ԉ����;�QPX�?2UE���(x1��EԦ���ác�p��������r<}�/��[����B6��@K*/9�����R�V,�܌��g*����z�8v�o,��U�@����=vy�|�a��JHEO���J�F�\��۠��Uq��$]��
&��L�.tmZ�;gd$Lr[�� g�>�A�
B�� ���3J���5�])�b����̾�:�����l��۩|6�����ޣ�v��#�|ԁ7��ѹd=��J�~�VC��~�֚��z�� �飈-k�=Ћ��@ s��k�yRj�Ĵ�.T�$�Ѳ_%Z�I�r%�H��[��A�E�P
/�<��]Zz@�7%��ޝ6����i;�F��I�7u����;A�E( ���+Hf������d9��@���Y����Ϣ�N�yp��O�@'������]�F���|��E@�(�[
��A9$(��Jy�����9�A�E�īY��f�7�s�F�T���p�
�?�0�d�α
ר�.���j�|N4�-����v�����5���d{&�f2�������D%��1P��c���@�&�pHk��V+r<������W�U�KGFm�܈���Vy-��iG�#�����M����]��>�jGS�]���ki"ӡ�l�T��փ�v�;��a��Dq��L�h�����ߒ���#�����4���(�� uʩ��D��)�]�0�Y�kY�:��[��ރ6D0�D�k/�&`X>��C�j�f�:h^sX�s�:����Nx�Fr���/K����,�*��1b�֒1�4�bl��=/�}�<41�����+�1�.�Z5 D��P��n��H~��maf�p9g>b�/�F~%��M�R�Z�C�`;��_����cC#�L�/8q�J��$�̠�/�~��b(�*��-�><�1���F�6kb�h0���	ml��~�R��ю�ZJ|%�;i�Iǉ%�._�8i������y�XW��?����=v9���rӉ:���:�Zr��$ݑ5�w�g�E̝�jR`)`�v���v�Lߧ��.n�g�j�C�g�[��φ�30ED%�lha$�|,�5%������|��(�2��Y��y�n��2�&�*z���P+ɂ��,0d,��t)���K)Dɮ�������ΰD2�8���0�|"���!WW*����岋F �����6����v��-�dք���Q�P������4=�I�t�|7��ՎL�-z?�{	 �1{2VM,�����l��oa�l�����a���ě(-ݚ̤�p8�*������s@��j�z����밁�G�S�C��g"lL�Π�XْD�c�;�i��Z���9������X&q�\�q*�4�K8�������X�gRO�ݞY��z˸�.�n"��|�jJ�莖8���y��'�'���|�C�i Q$�C�OKn���ܱ�.TK{��uVm3Ɗb_�S�ɇ^�L�L���V�<�ʪa��c�	��͸�LU�^�_E�l\��/����7m%����&'�/�^�{����B���̪Pԏ���T�!��綔���6O����s���R��?Hg��<��Fl�B5+�ө�Q2Uh��]����5�E�\ב�`�^�5}��m�΀-}����o[��w��l�[�ުU�-F��N��������#�Tb��&�1��%u������K(�����d)CL[�M� 9�!��"Qo��.E�\&)Lv���
���ի�����Y��=!�cV�z����b['�_)ˮ��.t��۲�Ӈvθ�C�7�'��"PQ�g�z�u���o6hi��F��,�
^T]]�ڞ#����X|�J+zbh& ����ʨ ��5M�D<�����ƶ���V�=��5�a�������c�;����eGZ�ȷipQ��K�j���?�J��Vp��I��ҤL�$��4��>5H�nnc�Tqu��c��0E���w(��C�ȒZ�A�\�d,0���}HvST?��b�#�g� I�*��e�	
 dHH�����L*���M� �=���x�7�`��TQN���_�82�q[��:���@Hd�)i2�35�pI��)����'Ǖ��%�~�v{IQ�@�yK��~x�R���=���D��y"�`K��'��4��;$�U���N�����J�AϪ���V��W��������|{45�x#�ӱ���Đ��vM8���='�/Z`>{W������Rl���Q��I�9��Y��M� �AuhMjG��`��X��Uå�5�c�� ><�pH��f�i]��O��$FYk��~W�T9��i>L��>���e��=�^;ւA�J��c�%`�N+oTY��-�����+��$\^��O)P��t��B4v%�^>��<�j�>t!"Nt�YF�/ϲ�/q}[[��|o_} �P(]�,�=R���|�3�Q�'�9��6��*н�?).����
֌�D�qԘ�Y
]r�x�z�:`V ڟ�ЗS�5�ߤl�oz�'�8������O�m�ED�Lb�P��m�l�U��33E�dǆ�Lԯ
�i���AF�Xm�0��TF+���A5�U�R���౵[�m��Ԅ#1��Ü
f��`V(�yQTNt�Q����YW�t�