��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL���m���C6%Z���[�$��]�IK�`�h�SyZ��:���|k&x��E?s��Ï�� �'lG��1�F45Կ(����Q��r�����L��R̕o�-:T�똛�u���o�	��M�͸��~�Ӧɯx��uxm��=�`HN1:ͅZ�{��Q�+2;���A��g�P�ȇ�}{�-Gs#hk���8�Ճ#��%j����x���G#����,8;�k�=蒃7bSF�f�슏���>��	�� =Sn���eZ���=��5�%o�
-f�W�fa����������ǼUTUK��T��4����\���^�l�-��a �0�v�h9#�F::z�}��$3��l�a��b(8�T3�S9�$	c��7ىRهwo?�ѽ�F]�{
���w�� ��I8.�AW[�����ʋ�AS
|��;����ۃ1���$Ґ�~���	����6�����:�?��B��Vt5���%�j?���A������-�)�	� ���݁�/t���SW�kn6�u^��J����u�;� ���V�l]�%����Tp�a����;��� 0'�L%,a�N��T�R^6���A���#�A�I���B��by솜*��<_��Cc!/J�/� �T_j9�����r&���Gs�u�$�G'y��J��Sr�z���,��`�yY��$�D�d��h�8)��v^i=�luT[��/�� �c=��!�c'��.�����1�/*~�3Q���fr5;�,.�H5�x]�� ��(k�l�&���'c4��9��k%F�f��E��|�d�xZo����Ĉ��=`����l7h=Q�V8U�`��k.қ*��ґJ��3 j5V�^ZB��w�e%����R��-Uc�?Z��g�S4������ �*�{�B���c&iK���ŭ�ʹ���8�.r���숯h.7�S�jy��}���?2nF��*c�q�4����`f��4��U�ED�g���ݚ��裙��\
��썡,R�������jۣ�Iz4ܶ�e=���2*7^�詮��3?R2dMT���(D���	P��]���3��]��H���S�刹'R�����r��6�C��bFCTwYim"�`���&�����2�n�rUE�R��ޟO�}�gW��,���C޵G��Wd�u+������#y��m��)ٔ����՞��Ͽ�>�������a�Y�1��ϱXh�/V��d-f�^�ˉ��?�s*wa*�QՋ��f��y�my���05���XtPSp��Uf�q|jc/�[�.�?��M[ٚ�t�9���ԑ	��i��h�ʸ�(�t���u^@��3D,{N�G��8�%'G��}�[���b�H6����RGu�����[d�d��=�zS������O��c!}o�4@I���o�4�>�s2c%���N{,�ڂ:)~��F%���"�`������;����_S������~��o�뉞���\a�p��h����>L2�R񔳚��U�}.o���*�v�{":O��{�P�mJ�?�m.U�Nu�TH�wcV�*�3�d�W��ԏM��.Y��o���:︧�%�j���b�"Y��Mi霉ݵ��q�v�?�1���X�yg��^�57��(��3��땘ˌ�/x���&�Q��J0f��>�*�4�)�\�F���AT��z�2%]=�G�axv��fݤ {L�3��S���K{�	TKh���t(�T�i�V[���th��
��s,wK�+����#jc�-YG.�}GO�Zo�
cl���^�ڰN�t��J���n� �c����Sk?fA=���UIR9���F9"����/#��������:�4D]��#�FX��Cp��n�q�ؕ�v�
��Ճ��e��O2��V/�u�C3�H$�X��2�y��cF�5W�	����H�#s�%`	t͜$r&�F��9 <�0�C���9Q����ςh��Sj�x3��E*��*��<�ޯA{P5�E���FZ�~Ʉ�k/�1U{�f����X��м�p��(�D���)?���Fa6N�q������qk2���lP�[{6�� ��OԍP�%������$s0��LOj@�f�L嫉 �T�w��*�R?<��h9�yAf��L�(N��ϲ�tu��Cuhb�^��J�ʕ�*uM�ЁZc]]�O���Hf�8����eR*xO��;���j�f=IT)��!�	Uq�.�~E^X�'LKX��8�]p��n'V�9c�iz.�br�r*-�i#���K���
��]��BYE*���{�ˠ%I�1rr<:�1ق��z���`=k�g
� �6�P�I>��Ԯw`��e]󭙸�b�����[��˜�����ڜB�6؍n.���!H�.�=�̐��W�n����|}��
vן-�&�5���9�tk|h�����X��D��P���>!q=�,/de,)p��b{U���1m�ف}�N��2
��GI1�pf�@�25�gW��I8j�� ��2>�)�,~�!�3�;]rʭT�D�R���Ӓ�2\vk��āN&2HYʩ!��������{N����o�K�����L\��*�a��%(�y`�AK�W���%�ܽ8���`2|�>٧_�X�%�4�M,R^2|HN{�X�Qt���]T<Ay&B%�o^�X�nsфn��TO|��T�.�4�R_0ٮ���O&�j�vshU��=g�� �ҥ��7bc_�ְ�?~��5/=�,�ؙi�������@�4��,�V��K(�{#�Y��FG�s�;�,�U|�"�M�nQ2�x�!]��}�ބ��y�J����y�p�l}�p�a	����܍v��NMѿy�HJ���&�ە)Y�ۗ�D�����?I�M�bo�ٓņ̾O}|z,l�]���2E �n�yH�������������".��֗�fb砞��V����G���ZZ����C�w@�c�a�s����>m"�!w��N�S�mgje�Ɇ��I��q�旴 �"})EvyY�t�TJ3�5r��
x�����t���ꕃQ�H�A�(�L�E�r#������v;�6���K���@�*MR�Is/�ϋF��<í�TI[O���
~(�ɧV��bD0Y�oĀ����[޴�n��ߡ��.��.��tY�a�~f`���=1�--�g���v�>��
DR�dJ$
�s5�_OS������&��9��)��}��b{��'��Yi�n]7�ק9���qդ�UQ�)�t�H
��n��Ȇ�&�G5���y�
Ђ�K �P���Y����.8<�'�M�f�~F�L�T��e{3�z��'���0����2�g�!�z̶�4��%<n�g�T[�W�.b��}�h��h�6�Q/�����苓ԱZ��A��E��%�����5�zl:��/�7l��Vxʠ���R�J�f�bt���ԃ�~�q0zB�ޏ�C�Ϊ���_�0��.& $޾r���0��A�S���Z�< T1�����������3�2A��9�&��!`�x
L�X�ڱ��g���f�*�_c�vc�Qz\�]dj���ɵX$}����8Ge�mp'��TL%��l�1�:���;������D�~��'؈'��s���N�sF��-�1瀃_���^Z�nT� ���$fV�K��L>pw�l:-m%������_	L%�yt\M`/Ш0³�p-�`�5�(s\��bR�>d�^��3���yZ�/�^q^ٔ��C���㾤�nj������|������L�[��Yw��/�6(�k�c{G[ģ?���	\}�������c1@�4�7_t �3"��� ]91�X�כ&�����?�xt�S��*K<M'�4�D�^��SM�8B&�֋�0K<�%*����Q���E�����0	����m?�Z�5����tD$���_蕅?�M� �rQ���㟡��ED�˴(M�	%��c�]���K�O[_X��n�e㕒��WS� ��J���:��Z�H>��i�8���5*ys�5���9ZDү���B/���6�%���->0�W2O{�N���"ߪ�$q������F���~�D!-�c4��t�R�yR���H���D|�,M�i��J����BQ= ��K����w��gRc�����n3)�Q
PA7G�����1�
��%
�KC�%���KпG��W����鹭7 zCG�g��/0�pA��S���)��5��%���m���f����隒��O÷�6�͐�^�L���z�J�A�j�uX ��\��:S�� ��3���$�:���5��J=P���5PO�H���C��;9�x�Wҕ���X7ku:�S�) �(�oj�� ]-�2.D�OC�8����N]��J�cc	0��I}l��2R�{���G��HeM��[N���}!���ϰ�����C◸x��'��[��z⿐��IPn�K:eHT4�I��
<����p;}���u�J��|Վ��{w���/�ﾳ��إ3n^��ٍGU2��1-�S�5�+螃J�r��I�]5�f�G�i��ZZ�g���-�\Ӟb����*i*Z�4A��8�v	�����a��@��'H�~�c�c%W�6�q�Q�Voʳ�G�v
h�pbp�0Յ�mW��ԧJM���>f:F��TSOl�������m�'g�Ҭ��!��3��
��;��]��T7�n$% �����pf��ƞ˴��c'��&�7(!���^�f�!!��a�}�v̖3����0H��wU����-���?�%�VO�U�2�څ�_O�N�t��3i����9��F��X��\F�]�~��M���� ly�Im�X�q�s�*00�<�������ÿ�>��|T�w�SF�cj�������?8��r��Vu��=!C��||��L=��ߛ�Mr�K��l�Ip�R���F�B6){�Ҝ�����cv��)M�
A���鿂�>��*r-��B̋I�gt2�T0b[T���`bV�����فW����]��L`45��\k�����W���k����#y�����*��m��� y�g�U�Nīcju�1�|i������mF�n~�����������	V�d�Qj`�uS,�v�Z��W���~�wf42o��+1Uv�J�5F�Y��B�B�����6G�KM�i|��7d�1u�S`�$���������͢S�lg�Gn�[�8�Z{ݬ"��$^(����An���꾺Y��m�0�����r����'�oD��?���UAH	tK�k�t�n���؉��@~�i�M��l>�@e�H����}b	�M��.Xm} �#��G��VL_�*m{���	�#"n3p��L���2����u�ۄ���]���`m�'��:r��׽��n�m�v��:ɧ� �W�"�\� �nG��Sa�X>�~ %�Њxp�2��V1F�4.�舚;>(��Ce��ܘ���˙CU�﨎YX�D��:�X��%ha��.��B�?N��������#"����=
��߇#�Kv�y�5���ݼ�2@�4�VI��~�� ��7�П��[�+�l�E�p6��s��[�^ѐ�9�ڏ/�׳{;}\�t�#��o�
��q��V� "�����cr�\6ha^���5/������ӈ�߀h3(5 Ө�\uo��m�2Sa�@uU� �e^gnT&��'���S4��Y��Z�S�NC`$Hnݠ�:y5�����Ԧ�R�B<1dw��}��k'�5�E�R�P` �n����մ%��pi� ��l�Ԃ
�:���cO��G��.�a��Ǡ0w���U�N}Sf�fA<��<�{�k�Ȣ6<m����\�G��n,��)b��� �M�;Y�D�o��b	a
��+�U��6�n���w�?�T��ٙƚWb�d>��		��J�PW��������$+�_=k��,��@;��[q�bY�;ezQ
V3U�c�x��5�۹��Ԕ��Cܼ��l9�.B������.�]�H7��
�)�9��F$O����d�_}���R�*{��h���j�u?S��	�W�