// system_qsys.v

// Generated using ACDS version 13.1 162 at 2019.04.26.16:21:55

`timescale 1 ps / 1 ps
module system_qsys (
		input  wire        clk_clk,          //       clk.clk
		input  wire        reset_reset_n,    //     reset.reset_n
		output wire        epcs_dclk,        //      epcs.dclk
		output wire        epcs_sce,         //          .sce
		output wire        epcs_sdo,         //          .sdo
		input  wire        epcs_data0,       //          .data0
		output wire [12:0] sdram_addr,       //     sdram.addr
		output wire [1:0]  sdram_ba,         //          .ba
		output wire        sdram_cas_n,      //          .cas_n
		output wire        sdram_cke,        //          .cke
		output wire        sdram_cs_n,       //          .cs_n
		inout  wire [15:0] sdram_dq,         //          .dq
		output wire [1:0]  sdram_dqm,        //          .dqm
		output wire        sdram_ras_n,      //          .ras_n
		output wire        sdram_we_n,       //          .we_n
		input  wire        can_tx_en_export, // can_tx_en.export
		input  wire        can_clk_i_clk,    // can_clk_i.clk
		input  wire        can_rt_rx,        //    can_rt.rx
		output wire        can_rt_tx,        //          .tx
		output wire        can_clk_o_clk,    // can_clk_o.clk
		output wire [5:0]  segled_sel,       //    segled.sel
		output wire [7:0]  segled_seg_led    //          .seg_led
	);

	wire  [31:0] mm_interconnect_0_segled_controller_avalon_slave_0_writedata; // mm_interconnect_0:segled_controller_avalon_slave_0_writedata -> segled_controller:avs_writedata
	wire   [1:0] mm_interconnect_0_segled_controller_avalon_slave_0_address;   // mm_interconnect_0:segled_controller_avalon_slave_0_address -> segled_controller:avs_address
	wire         mm_interconnect_0_segled_controller_avalon_slave_0_write;     // mm_interconnect_0:segled_controller_avalon_slave_0_write -> segled_controller:avs_write
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;           // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;             // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;          // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire         mm_interconnect_0_epcs_epcs_control_port_write;               // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire         mm_interconnect_0_epcs_epcs_control_port_read;                // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;            // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire         nios2_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [25:0] nios2_instruction_master_address;                             // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                            // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                       // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;        // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;          // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;            // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;              // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;               // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;           // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;        // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;         // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_can_controller_avalon_slave_waitrequest;    // can_controller:avs_waitrequest_n -> mm_interconnect_0:can_controller_avalon_slave_waitrequest
	wire   [7:0] mm_interconnect_0_can_controller_avalon_slave_writedata;      // mm_interconnect_0:can_controller_avalon_slave_writedata -> can_controller:avs_writedata
	wire   [7:0] mm_interconnect_0_can_controller_avalon_slave_address;        // mm_interconnect_0:can_controller_avalon_slave_address -> can_controller:avs_address
	wire         mm_interconnect_0_can_controller_avalon_slave_chipselect;     // mm_interconnect_0:can_controller_avalon_slave_chipselect -> can_controller:avs_chipselect
	wire         mm_interconnect_0_can_controller_avalon_slave_write;          // mm_interconnect_0:can_controller_avalon_slave_write -> can_controller:avs_write
	wire         mm_interconnect_0_can_controller_avalon_slave_read;           // mm_interconnect_0:can_controller_avalon_slave_read -> can_controller:avs_read
	wire   [7:0] mm_interconnect_0_can_controller_avalon_slave_readdata;       // can_controller:avs_readdata -> mm_interconnect_0:can_controller_avalon_slave_readdata
	wire         nios2_data_master_waitrequest;                                // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                  // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [25:0] nios2_data_master_address;                                    // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                      // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                       // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                   // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                                // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire         nios2_data_master_readdatavalid;                              // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                                 // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire   [1:0] mm_interconnect_0_can_tx_en_s1_address;                       // mm_interconnect_0:can_tx_en_s1_address -> can_tx_en:address
	wire  [31:0] mm_interconnect_0_can_tx_en_s1_readdata;                      // can_tx_en:readdata -> mm_interconnect_0:can_tx_en_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                       // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                         // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                           // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                        // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                             // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                              // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                          // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                     // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                        // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         irq_mapper_receiver0_irq;                                     // epcs:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // can_controller:can_irq_n -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_d_irq_irq;                                              // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [can_controller:can_reset, can_controller:rsi_reset, can_tx_en:reset_n, epcs:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, nios2:reset_n, rst_translator:in_reset, sdram:reset_n, segled_controller:rst_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [epcs:reset_req, nios2:reset_req, rst_translator:reset_req_in]
	wire         nios2_jtag_debug_module_reset_reset;                          // nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	system_qsys_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	system_qsys_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	system_qsys_epcs epcs (
		.clk           (clk_clk),                                             //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                  //                  .reset_req
		.address       (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver0_irq),                            //               irq.irq
		.dclk          (epcs_dclk),                                           //          external.export
		.sce           (epcs_sce),                                            //                  .export
		.sdo           (epcs_sdo),                                            //                  .export
		.data0         (epcs_data0)                                           //                  .export
	);

	system_qsys_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	system_qsys_can_tx_en can_tx_en (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_can_tx_en_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_can_tx_en_s1_readdata), //                    .readdata
		.in_port  (can_tx_en_export)                         // external_connection.export
	);

	can_controller can_controller (
		.csi_clk           (clk_clk),                                                   //        clock.clk
		.rsi_reset         (rst_controller_reset_out_reset),                            //        reset.reset
		.avs_address       (mm_interconnect_0_can_controller_avalon_slave_address),     // avalon_slave.address
		.avs_chipselect    (mm_interconnect_0_can_controller_avalon_slave_chipselect),  //             .chipselect
		.avs_write         (mm_interconnect_0_can_controller_avalon_slave_write),       //             .write
		.avs_read          (mm_interconnect_0_can_controller_avalon_slave_read),        //             .read
		.avs_writedata     (mm_interconnect_0_can_controller_avalon_slave_writedata),   //             .writedata
		.avs_readdata      (mm_interconnect_0_can_controller_avalon_slave_readdata),    //             .readdata
		.avs_waitrequest_n (mm_interconnect_0_can_controller_avalon_slave_waitrequest), //             .waitrequest_n
		.can_clk           (can_clk_i_clk),                                             //    can_clk_i.clk
		.can_reset         (rst_controller_reset_out_reset),                            //      can_rst.reset
		.can_rx            (can_rt_rx),                                                 //       can_rt.export
		.can_tx            (can_rt_tx),                                                 //             .export
		.can_irq_n         (irq_mapper_receiver2_irq),                                  //    can_irq_n.irq_n
		.can_clkout        (can_clk_o_clk)                                              //    can_clk_o.clk
	);

	segled_controller segled_controller (
		.clk           (clk_clk),                                                      //          clock.clk
		.avs_write     (mm_interconnect_0_segled_controller_avalon_slave_0_write),     // avalon_slave_0.write
		.avs_writedata (mm_interconnect_0_segled_controller_avalon_slave_0_writedata), //               .writedata
		.avs_address   (mm_interconnect_0_segled_controller_avalon_slave_0_address),   //               .address
		.rst_n         (~rst_controller_reset_out_reset),                              //     reset_sink.reset_n
		.sel           (segled_sel),                                                   //    conduit_end.export
		.seg_led       (segled_seg_led)                                                //               .export
	);

	system_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                (clk_clk),                                                      //                             clk_clk.clk
		.nios2_reset_n_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                               // nios2_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                  (nios2_data_master_address),                                    //                   nios2_data_master.address
		.nios2_data_master_waitrequest              (nios2_data_master_waitrequest),                                //                                    .waitrequest
		.nios2_data_master_byteenable               (nios2_data_master_byteenable),                                 //                                    .byteenable
		.nios2_data_master_read                     (nios2_data_master_read),                                       //                                    .read
		.nios2_data_master_readdata                 (nios2_data_master_readdata),                                   //                                    .readdata
		.nios2_data_master_readdatavalid            (nios2_data_master_readdatavalid),                              //                                    .readdatavalid
		.nios2_data_master_write                    (nios2_data_master_write),                                      //                                    .write
		.nios2_data_master_writedata                (nios2_data_master_writedata),                                  //                                    .writedata
		.nios2_data_master_debugaccess              (nios2_data_master_debugaccess),                                //                                    .debugaccess
		.nios2_instruction_master_address           (nios2_instruction_master_address),                             //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest       (nios2_instruction_master_waitrequest),                         //                                    .waitrequest
		.nios2_instruction_master_read              (nios2_instruction_master_read),                                //                                    .read
		.nios2_instruction_master_readdata          (nios2_instruction_master_readdata),                            //                                    .readdata
		.nios2_instruction_master_readdatavalid     (nios2_instruction_master_readdatavalid),                       //                                    .readdatavalid
		.can_controller_avalon_slave_address        (mm_interconnect_0_can_controller_avalon_slave_address),        //         can_controller_avalon_slave.address
		.can_controller_avalon_slave_write          (mm_interconnect_0_can_controller_avalon_slave_write),          //                                    .write
		.can_controller_avalon_slave_read           (mm_interconnect_0_can_controller_avalon_slave_read),           //                                    .read
		.can_controller_avalon_slave_readdata       (mm_interconnect_0_can_controller_avalon_slave_readdata),       //                                    .readdata
		.can_controller_avalon_slave_writedata      (mm_interconnect_0_can_controller_avalon_slave_writedata),      //                                    .writedata
		.can_controller_avalon_slave_waitrequest    (~mm_interconnect_0_can_controller_avalon_slave_waitrequest),   //                                    .waitrequest
		.can_controller_avalon_slave_chipselect     (mm_interconnect_0_can_controller_avalon_slave_chipselect),     //                                    .chipselect
		.can_tx_en_s1_address                       (mm_interconnect_0_can_tx_en_s1_address),                       //                        can_tx_en_s1.address
		.can_tx_en_s1_readdata                      (mm_interconnect_0_can_tx_en_s1_readdata),                      //                                    .readdata
		.epcs_epcs_control_port_address             (mm_interconnect_0_epcs_epcs_control_port_address),             //              epcs_epcs_control_port.address
		.epcs_epcs_control_port_write               (mm_interconnect_0_epcs_epcs_control_port_write),               //                                    .write
		.epcs_epcs_control_port_read                (mm_interconnect_0_epcs_epcs_control_port_read),                //                                    .read
		.epcs_epcs_control_port_readdata            (mm_interconnect_0_epcs_epcs_control_port_readdata),            //                                    .readdata
		.epcs_epcs_control_port_writedata           (mm_interconnect_0_epcs_epcs_control_port_writedata),           //                                    .writedata
		.epcs_epcs_control_port_chipselect          (mm_interconnect_0_epcs_epcs_control_port_chipselect),          //                                    .chipselect
		.jtag_uart_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                    .write
		.jtag_uart_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                    .read
		.jtag_uart_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                    .chipselect
		.nios2_jtag_debug_module_address            (mm_interconnect_0_nios2_jtag_debug_module_address),            //             nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write              (mm_interconnect_0_nios2_jtag_debug_module_write),              //                                    .write
		.nios2_jtag_debug_module_read               (mm_interconnect_0_nios2_jtag_debug_module_read),               //                                    .read
		.nios2_jtag_debug_module_readdata           (mm_interconnect_0_nios2_jtag_debug_module_readdata),           //                                    .readdata
		.nios2_jtag_debug_module_writedata          (mm_interconnect_0_nios2_jtag_debug_module_writedata),          //                                    .writedata
		.nios2_jtag_debug_module_byteenable         (mm_interconnect_0_nios2_jtag_debug_module_byteenable),         //                                    .byteenable
		.nios2_jtag_debug_module_waitrequest        (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),        //                                    .waitrequest
		.nios2_jtag_debug_module_debugaccess        (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),        //                                    .debugaccess
		.sdram_s1_address                           (mm_interconnect_0_sdram_s1_address),                           //                            sdram_s1.address
		.sdram_s1_write                             (mm_interconnect_0_sdram_s1_write),                             //                                    .write
		.sdram_s1_read                              (mm_interconnect_0_sdram_s1_read),                              //                                    .read
		.sdram_s1_readdata                          (mm_interconnect_0_sdram_s1_readdata),                          //                                    .readdata
		.sdram_s1_writedata                         (mm_interconnect_0_sdram_s1_writedata),                         //                                    .writedata
		.sdram_s1_byteenable                        (mm_interconnect_0_sdram_s1_byteenable),                        //                                    .byteenable
		.sdram_s1_readdatavalid                     (mm_interconnect_0_sdram_s1_readdatavalid),                     //                                    .readdatavalid
		.sdram_s1_waitrequest                       (mm_interconnect_0_sdram_s1_waitrequest),                       //                                    .waitrequest
		.sdram_s1_chipselect                        (mm_interconnect_0_sdram_s1_chipselect),                        //                                    .chipselect
		.segled_controller_avalon_slave_0_address   (mm_interconnect_0_segled_controller_avalon_slave_0_address),   //    segled_controller_avalon_slave_0.address
		.segled_controller_avalon_slave_0_write     (mm_interconnect_0_segled_controller_avalon_slave_0_write),     //                                    .write
		.segled_controller_avalon_slave_0_writedata (mm_interconnect_0_segled_controller_avalon_slave_0_writedata)  //                                    .writedata
	);

	system_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (~irq_mapper_receiver2_irq),      // receiver2.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
