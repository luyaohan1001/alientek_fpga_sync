��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ���$��`��:*Do��@f^)���3��de�3EZ�i���@UU��j×��)�?��Զh�&�����y�����������^㯘�L���[Vz��͟���B�"����І��Oo#�~�GDJK��ص!�"p�\� ���N�A���j�vbJX��8�
�D�� ���I��Qx�X����"n�e�x�`#t�qO��9K's��df��]�]���NoGʭ�t&wedc$+��%+e#Z����4���i:
�n�����mLJOW�Z@kx@���G�]����D�,?�o�]1�yuN�)v�H�	�>Je��@�_
=5�^9��p?���rی�E�޺��.��1ƓTPl�����2T����
Vy5�'��Os��|UB�Ssl%n���uYjh㕼�$\���\�/rD���8����K�[^b\Iy��=��":)zs:%������:�T8��%g��zk4f����-����=VWm-��QV���=���|"݉>v%nܹ�>��,����x����v���P�����拵�\e߱+�����RJ��hjо$������PC�h�)ٜ��>k��*]�T�H\�\?LS�yFG�H�ؿ�B���H��O'������&j��C��j;����SMG���Ȅ�����;`�Z�h��3�K�b�ؠ�3	<���hBS�U�թ�� <���A�J��	���"�b@���l�O6��0�l:������P'���,�I���4��y�Ih&7����g{��B��Pzq�}H���6ת�ӃX�wF,�(�Ê��~�77�a�~VW��`f���Ga6�U8d��d���@<�A���
_jVߥ����AI5���a�L���1��o{0�w5ۧ���5k��錑L�-���g����:�W������(&�$O��&?+�3�"Į�!p�˺A/w�n��>�H��� "������m��v���Wd�h*F��J�Vȍा����=	jqU M,�0C�?!�|�1�b�sO��K@���ͩ9�M:�����+�ۂ�e9m�e��[U����9W��=/�c�+�P�,�7)̏�pG�[���ko��K3S�:Y\+-0�
��9mƆ��n�@�f�l����t�I`
���M��z��	���t�Z���U�d�`��\ku.O�����Qڪ�jW`�U�Lw���z�M&P@������Y&�k�{�$u��k�&�gq�;�u%�f�ՊX`F���W�x�r��W�f\C�4ER��isjm9����3ō�T �@���&/��+Nf�TK��"�ۀ�hf#g�q�%<ܒ%��~�t"�>jtjޛL���K������Ӈ�����^�#
�&��M'xD���JO�̩R&	#�g��I�N�퉗���?h5ml�CZPں��]7\�|sx�w�{���㰸�4nGi��Et��D�ަk%�s��Pe%��z���H=���85'?dw�Z����#�:���F/MO�?���9>�>�r�:��݂��L�X� ����RH0E|�F�hܨb*�?�y4��x�	^���뽃��(<�o0�j"X�?�N��̯ͭ��Q_���n�8z3��nL~�vN�0���(�:<��t�% ŷ���jV�-Œ�4+$�G
ٞ*ۛ`
^>�V�n�}��0:#�^&Z���a_tH��Jڣb�U��!�M��MwcF����("��>��J5���n��q��g#�c��<�$�Զ,����=�F2���}�k�]1B�GN�?���f�4���~Od=ܚ�l��M[ˇ<�(����8��s�s�K�9췈}�$��vUs{N������LA��%^���TG��^g/���B�0�(�n@�XW"���sq��J__e�z`R; ���"H
�����ř�����S#@,��M_�3�wf8�T
JY�s�/�\XA�h�V���@s7�L�50��v �K�Z��n��~�ߕ��ޒ�av�2����[�IMP�-3��	|KԨ���������'Q��D}�������)���I������'�=�*��������Z�7g�����^�G�U��_�Ȣ�ݟlr*�E<n7}���m���Y�1��˫��8e!��sA�����1�D��|��I�4���:��+��5d��1{�i��0�O�>��a����֡�{�}�O���vw(�O}�����3��9�(�o%|� �6l�|L7}����s-&b�H�!m���1�:�GJ��N��cw�k:m^�\fh1G��� �ˍ"�j�w����3mH�	��
��C����ގ����Ճ-P� m1:�|p�q� .�V� m@���#�c�A�)�O\���\F�q~X�{b"9L�x[0P9�.&_�Y;Qŷ#�45r���Q{ٽ�=p5d{�b�'V���NH�Q�)/Ʈ�;�u��R�r�����տq6�+�)}^�4��-���o�ݱp���$؁�}������i����(@�A�~���1���G�ZѫT�n�ID_f����ø�����^G�����7
��&68��F�epk��|��2iF��5yAtJ�����gI�Mg*�Qƈ��r�X�/�@	*,{朠�d"3�R�_�s�Zm�z���Q�5_���������N���M�Rw�͸	aE�����j˜�8�T���P�Pn<=�b���1���qo�}��
����d�H��:C��q4qB'S흷�n�	,9��[��q1�D�+y��4�K�*|��dX�������G-��
qHfkBO�</fi���ͼ�kBƚ�`���#U?�{�;��|� E�My�b���+O���!��#8f*�M�1+֮}�NE�w=��vȷ�I���;*�E!_�o�]�|�Lp�p���E�"
�ߓ����խ�#����:v�ߍR�����g�I�H/��Yru}1����\��8�� �T�Z	d ��sQEb����ֵ���K�<��eB7(�D�ʳ� �p�#�� ���"^ۣ�L�r��t�QJ}l	0 �J���h~J��\OG����88��ψ6Y�
��9�S�Q���PĎ�47`s���]�(4��c�8/���&$�6Ԍg�����t�;�{ d�-_���_�)BXj!��'R�h9� :'-FU�`d����
q�.-�/	�ة��T>�h�"}?�0�u�'��xn�<^��3U�h� Y�mSod{\�p80�����]̓�������w+G��l�Y�%���{�8��'bԈ���3S�g��
uzB��	�v���]�Ȃܲ�Y�uަ6���� ���=�8WcAL�8�#����0�@	�����h��m��<)�Ω�`�0QJ'Rk���l���#�m�L\\�2]��� 8�V��p��z1UQ�A/��=� �`��X{2����7����C�����&D�&���a�+������h�,qbJ�W����(4%�)�W$�ܑK�h�O�֬ljq�1��Is(
��{��$;�*J'�m�B�ӊpp�F��q�����^����	���H��l+�����p@���t����H�����}pl�mک#&X'��]���r`}���`-��8ry^��޻�� ��(�M�w@��2ǕYk9ȧ]"�1j����O3:M+H�% ¨� ���nE�+�Bge�)�t��!Nx�
���� uK%5�IJDWhF�e'�R�����q.̽��'�%(x�à$������,V㽖����s�G�j�A�^�
ɒ)���%�욳�frͨ-� !���r�[��!�DZ�R6s>a]c��H8O�ӈ꣇��"͊��A. ��ת���I�Ǵ�O��6�a���� Xt�V�E�E�_�����w�/Ab�x���*�Z������JSǨZV�
��kݦW7VqsK�?��\�y| �˜�8e�C�~�$�����k��sS��/�1�W#/�|�`��80���R�D4�nQ��ȹM���b4��FX��Bl,�&"*<0�cC�؉ƍw�- rh�!>?|3$O�E�F�t��UI���K�_@�Q�Y�)��2ǐ=oֶ����TBc� x�i��F��t�נl�\�o$uL�)����8蔌W��+�� �gC-&n���r�����Z+ǵ����.G��b��w"	���"k��OdKl�%��oڣ
3Ma�y����Tڻz��v�K@[d4<[�_�QQ�{�#�'��W�
�F�����o�q����Rgvg��\�LV��d�J��]\���A0�@WW������9.L����]rڊFb�`�w�c�,�����jD���Ѫ�\P�;�\��L��` ��o$�a?�'pv��	S����b_t{�&�0��6��A�؅��M4t��X�w>����]�;;eᨵi5�l.RY���M 1�܃]D���j��W�k�����?j|M���_˳�uăy�A�<��ٴ��TA1�+��n�9�P{uK��%�$��P3�����'�Z����(�l�RX�%�9��'&�{���&L��j���� Z�V�uoPE|m�������8����~�ޢiF��GЬ�2��Uâ�v�֟��Y�1Wޑw
?����L�����X8���T��������xQ�U���븟�a�D���2{�[�J78��y� |�k��~8���D�f��e��r�"Q��v�� �� k)Yo�W5��(c�4v4<�p[�Q��z����	e��/��9�� u�4|���Ug�rVe�d �g[~:��8�n���h '����n*F���~f�NP?�!k����筽�#eUR�״� u�j8̄w�/�|<Z!�+�J*4�DdT��ِ�z,[��������x<�ϠdFD���C"�eй�;�u
�^JnIbg����M�ƬX�7�����Q��OOE���0뻌�#+�".PA��R��PN�6�Z#m߆:� ���\����>�̿��l8����n4�̿���")��YL�!�i���?Qzz�z^*��yQ��o>�5��G��|Td(��P]��7ő۸2� N,��k��x�s��e����;t�S�izmu ��]��x�^���l�nc��v�޺��/�&�\��n�{hJ�b��z����s;Yk1y#�S
e�7T����S�p�F�Ҿ�5�P�b�eu�a(t�ͦ�{�=�,X >�B�aE2T�j��ӻ��V_�+�D��m�lk�=/6-}��R��,���1��[LT��3�{n���m�%Ij,yxm��Ń�;�n��'nI+��"����-+4�����m�#W˰��Ǘ�E���e��;�>Sjt3��<Wh�#��ԶO�		0�{ɽt�W��~����P����$ڻ�*NM��{��ei��N|咕&n�N�pH�&*��j�@���&�D�S����vCG��<��s]F��R�N��OPՙC�Z'L8,�������?��&���Z�A������ń�ˬ�&�=��%Í��{m�)"y�����,��S��
��;d׌�3IW(�t1��]��.��*iD.b��+�*�A���=�b�:'����@d4��L���.�Z��65�6�[����[F�]Ð|aEe@n�S� k���ǐ)���<�b���(��+�m5���j��q �c6QA�?h[.�
�#�^Pw6��'F�,�S����\�3�LO��A��p��ע#���pi�H�m]U�<��oʮ�?^E�w0�O��c6�+�b�����ĈԀbm��N�j�䌳�<���������,��H SD�w�8���5��^b��~Aa�xo�t�`������k`l3K�1t�xj��u�	�AZ�z��=AHb{؞fy�8$$�77�ި��ꗳ��;%�z&7FA8���O,�ƑFf��۰5���,��,AX�=�;mȑ&�t'*=����ε�Yrۥ��t=�J#�%�5~����p���Q��_�K�L�l��1��AFK�&M�9sFL���:�c�"|�Să����BA����s�H��_�V��۷1�+��,���8}P�<"o�=�|,ށ��ZV��y���������1��@]�`Ui�&�����W�]��[�lYԬ�)��e�<����։�K�wb��9HB9����֭�{����r���o�������p���sn��n	 h�i��~�3�kJ�?�QR��73�3�x5��C��Y�Z�=�q�����mo�a�K6�5@*!O�HE%%+\ė��o��d!��Υ���8��=%8�H�|����ի=�S��������h`����{!�ݤ׸�vg�� ���2�m�  �"(�`�EҌ�T��lM��~c��C��a����Y�cw+Dt��*�+�[t�犳O�9M��g'L��鏎;?���*J�
�f��z�R(d�;��rH��j�Fx-��Ɩ���%i	m ����M;>j�C�~�Ȕer�ǸW`�Qj0�yK˰� ��>u��������di�wjp��F����;�4#����n��o=��CZ?->���U����9dL[�naXaw�ݒdl�+�������5��Ѱ�d������Hr;q���:$�xW��
�w�U�&�98��|�n�ش�#��n� ��ŀ|��v�d
�^�{�9�(XZ�K�$�ˀh�������w�(:0)|��P	�$u���0��¢�H3�jD�u�RS�h�0��AU �x&U�n�r�\`[��3�]YOp��g���>\��L_*O��n�f�>W�qx�ߺ�Р�9Ӓ��5n��5T�������t|S*��5&�rU͛*Ji��D`t�y"����޵�q`���:N2�E0���s>�6?�*�%�7��$c��ٙ�~ݳNpp�#ʹ�d�q�tE�e�A<B��=������m$� PaN2����F�qu��`��=j_S[��
�JF��凗���R��<j`�Pl��u���6��TW8�>�Z�����ml�`��-T��3��eo"���xc)Q�cw��7b�Q�����wϴn|�+��v*6�����j�l�5�N� .k���F����y>�F�;����N �0$�V�[H_v�M��EB��쥚E���WA�-1.���D���jY�(f�͊�y_�
�(���#M�&R�l�������;>�ʬ'u��LC'��R=�p2"��8�i�vt��)C;������Sɩ\1��,�Q�3
�P���=m"bzV������?�i����y�הñ����w
#��[]�ѥ*W �2�~"\�<��06_�����?i�z��$�`l�͵z��%��k��mXy�ò�D��N�,��ۮ��}�E����-�_�G6Tm*ã��pN��^��m�H 2��E7&_B �͎0e���EJ�y�;:ewX*��T$��̽T�`��'G�6|�H��� �Avc�Uo��"�u�w�X�v���&��őR!�	�ԧ�>+�K�wdv{ ToGF�R��QH���č<��Ť�ؓ��ϗ{�;g�9��fc��Y'��D��7�����\h�Ru#U���z?�N�ڗ�|5P��Q 5�&��Y6/е&�]<䑮��L�;�l��'���"�*&ac��i}�Hl�k�\�6��J>}nba���j��Y�ܫt,H��:��ؕ��MI�;��e����
3P�1O���7�߸/!���^�x��g]O��U� �g�M�1��VQ2crs@A{='�EP�����G��ԕ���;�����R�/���]�����`9#]gg����\��P�u�}�R�	,B2㺈�Ym��!��X�c��۝�t���ZMUO�!�������΃w�����c�]qH&`Ѷ���z,`%�e����"�//<�}T�\V�'�wG�~��޶�}�}�Q�u�uf�ݟRB\M���:y��(+y�}�0`�d6-C�q��X��#r�%1�=��񧭍Z�9��?7t���K�����ǥ�c��z%f�o����R��;�V80���`�^���zP�
%��
��9{qM��/��u����c�A+�����⵭K��7U���D�7��dN0D���}p�`��M��[WX�`�"^���9�=����r%H]~�m����[���IlV�쀚����69Ō�rZ�ˋ�nn���NO����]\��[D
�&�+$����A[^EO	�m<�78�'�2�}b2���ك�X�X�oN�%p\����\���WM|�����K�O�"���&Vu�h������M���ʚ�(`g\�AZ��/�����<�>X�xVf�|�]�:b�H��H��8n*�^3�4�U�F�x��W�IH�'�ne)�[�)dG]�V�*ܧM�K�	c��K�sc�6�׿҈
�G�H~>j���w֗�<:M��aJ���'�X�8�e�)*ݚ����M�8S����}�u�Q��1�#'Mz*��m
dLf�c<t��I,M�;n|,6D0�3�{7�Ի�X/[O������k0�"b�����k���Ʈ�� �����@�i�B?+�y�gp�B�����<��9O%s�`���(�srR�<ZDBr�4���EDIo4['�f�����`�?:E͙�d��T���i�2�KJ߳`
v56l`:n�&��7~���E�xK�AaAx���`#z��8o��PTc�i|�����^Su�K̱ctxy�:ԓЬ]T���LL�K��Z�f��_��V����ǋ&@���t��c�M3-�K���vS@(��RZ%����#D%�����,5��t@lA�{�md�9����Q��j�	����H�sk3*>�Ӫ��aT<p���SL�Q�hV����*�Ģҝ���,*'�#-����K�S��]�Ԧp�7F�߇1��,���РH ��ceV�;�}�P]�u4�~g�ӫ�i0�wi�?�ᭂ�e�y#`�l��aR��4'��I�G�ڹ��Oހ��^?��8TK��](;��|�����Q�]�}f�,�[Q)%<LH)H�ޕ´�6�Q�ݧ,R�ho?*8���8@�J���n��71ː���1;�G���{bp��Ά�����z�q L��5����0X�;��%�b�2/�iW�_F=���ƈ�#ުG&Î��.o���a�@��Γe��1re�4����L���p����l����P:�DӞ#~M�m�䪊�3�Z[�=("⭡H�V�龭c�>��Ao;�LQ�̢�C��K`�1�Ȩ�e�n��ioJsZ
J6M�dR�R�`��$r��zO:�?�VvsԈ���,��nx��h=�ǫ�N�rK%"�9�8rM�Y`}z%:�5A���4녂��13�ba�R[|K+�i��l�� �Q�L"E]dn[���A�?֖6�OƁñ�V�(+�q;S7�Y��z����)���2F�x�ř����g�T=��7�;��_B=��d���Z���Z���7��zm
��z@�(	>cE�����)�qa6T[-�F�J��, =dy����=Z�f�yư��2j	��cLvd۞���Tz��O5����Ul��� ��s.S�?�ο)�͏�ك<	�̓�<�߶��9�KP�s�u9��I�1P��_L�����c{l��7K;�@L��H�Z��E�;�\vt�r�	�i1I%���OC�H�R�Uc/>���;(e����WZ�u�<�(#W��;��3 �黺�U��D�ԡ<�	i;$T֓Dx�=3�{�p���q:���aK~�x�� Q�w�Q�R����"�4#3�u�>̢�^�ă��`�Z�4�	pw�"!�g)�e~4�v�>Ǎ��qc����c �[�D�����e��dA$}�:`{f�p���v�>4l:�!�4`NV(�)���a���i�-�.(
ų�4:��q��J��Nќ�@�˯g��T0�.̄L=��@g7I��,΃/���)1Q�ϥۜ�jw�UNP��X5�\�X�i�I]���D<Z"�~i�1X���FzB�!���W���v��L���h�3&%�փ�gD�u�(J��w�g��v#�t��*�؜Sه�G�������هR�Ҿ׊\�(t.Mc~�) i0�:}�۹ 4�0p'��E�-�9�%�`#�hw���ެ�˓�z��^��/�8R�\APn��ҷ�� q�g�j�#��t8�c��¾�np��da�r���d�|
����27>C�Ll����7>��NJ�ʡ7����R�h�<�ui��+V�AO7#s&?f���'[��C\�?T/����?�PH���p�D/$YL*�p^��L�'*'A�)��.�-�0PJǟz/iIb�y��< ��:U��P/��(��ގ��t�W�n]�)&HqOB��=^2z7�KU����oњ����2.3��Z����2Ձ�Ix�/o6E��i��"ϑX�v�3��NE�'��x��'=����� LT��$'	�o!����Q��͉������ז�<�/�Z���qw�4!6g��4�z��d)	W˲\o����H��[�C�q�ښ���j���U��9]l�����\R���M�5Hr�� f��c�R������(��!�v����32�V�jE�J%6Ԥ;�W�0t�� s0����q8�'oΌ@�8s�0�v�]���'u��9�30҆�Q�(r-!<u��/�-��W��P�a���-E�%ԑpIV�{�d����0$�������BU,�k�\ؠ~��V�Zi�bS�{�p�|3�'� q��Ư�O�i��d�]��>�H���e`p�V��u�?�	����tJh����2]WF�d�.���)rpW�Ľ���$d��`�0�c�-ZhQ�8T��/�1�1!�E�*!�GŒ���}��VVX}� )�	x���)��?�*��k$��Ǣˁ���XB�6�ݕ_f���0܊+<E������0ʷ'_������,d 4}~�MZC�+� Y��O���q}��Hv���]��Lm&~j�r:�rUH�[L�s����7���!�dŅE�wN�♘1�I�c���/bD�CX��TP��c3N��d[OA�+�n�]��*C)ð��Y�O����;=@����Ŵ���^ҩ�:�+��
������ׂ�:��O���6�D��3wL+O���0�n��__d����\ꋫ��Հ���ê����Kp*k�yZ��;�X�7z(ч��:��sя-��I�|C��WN�Q3���^\fs$}J��h���V�.��~Gh7 �p6 ��S��?
B���erj�0ga���!�i�b^|���j�%ߣW_�b���7v�]���ˈ�HeT$�5^ �ᥘ���p1.Mb�g�R�(�hҿ�=�q�}�9l_ٷ/'߭�f{Xt���'g��b���s�1�Q��q8ڍo5���|�E�_~Eu��������N&G ~��.��;dᅇ��B<��P�%�f�/.�����_SG��p�6�X^�����%�.�r%����xVL�_y����Ι���	��g����l���'�ĸ�vF�&��1���J�{��E�àl�� T�u&+��jX.蟻����~7QD�r�:�{CҨ��̈���z�����S29�2�h��m,	�u�ǀp��;�tX�'5Zh��tx����� Ү��򒠀��D��g����y���.Ϳw��Z��zG��X��t%��#8�%�@�w$JV�F�E}N�=C��l�G���Nuv�H�)�,s�3�ѻrD_S쯰��f85�'��d�x	J�L��E�{��9`�I-=,� �i,�.r�-�CȣW��E��-�_6��Z����=�O#�]��މB��5�E�`5����N@�G�C�RW�� V/J�L��u��e����A��H���27� �I�yv�`�`B�]Z��)i��3������9V�JQ	z#� 1Sd�u�|TP��49�?T��6ϝ�e�)�[w]]oj, ��y M��I7F�+�b��@�b��$}=�F��FE~e����s��X��d���a�#,n�6��_=���U�2��kX�9}p�a�)�`�ť����,u���+ѩ�q�4"2��5=�w�!���+k�fW�ɝ��zr���DLр��NB0�V
O�+y��?1� �Ł�������P�(��<����vV(8?R��Ij�(�j樣r$��is��Ld����\v���,���5
.���[�8r���a �Z�b���Ws;���j��s�����JO��y��p(KgU�̩�E!��fLB��t,��O^>X�F�*�	W�B��ŗ?�۔��������GW�9�{H�wQ��Ĵ�U��Df.�����z��O$�|4��S�,���B�p�Y��T�~bK��:"7р}3���p͖�::VǍn�M�u���}��oݺ���/��ǈ%�Z����6�ܻ�N<5�_=f��"���҃�O��ϧ
����8�5 朶f����
���q=E�1�c��f�5�b�iVﲘ���[&{ �L�Ry�����x��+E*�	a�쪉���L�*�j���xd�׏��` 펎��M.N�$w_��3�=_���
��Y�X�5���G^I�삫�òXp�M lۏ��_�&iP	zs�?���|�ϙQv�
�
 "�=��L���P6�:o�F'���2#�g��wF�2	8��@?,qj��LrA �1�g��LrL�S㪰�5 ��Ea�f�*����(�b�>�1�G�Cr.�إ�������������@�NǧS��a�b��e�u�bM�������N
x/�^,򪘟0����D2<,Mܻ�ܨԋ��n,,����ܣ��"��wI+�!��?�d���[5:�ΌR�B�����94h�@�!rr�����t��� a�R�0~�M!�0��;y�K�U-7������h�"dF������z0 {?�t���������������l�ʟq�d]|�2J��J�i0�Gڼ\�ѣ>�a�IJ�"����PfGP���e�H7�Bҙ]nX��Io�p�S�[� ��$�OX���ż.�&Z@�}�ၶh�����M��z�Թ���<������Ӏ}"����%�\�8�-;��EI�J�\u�/a{VO��>��p�4��{��B�
�,���35����U&�� ����N7�b�D�5fhA�E&|��߉ zUU���O��r((�D�Q{�ҥM^+-�.fJ|q��*�,����ċ+==�Zטz��_����aH΢G��ϋW���d_�ω��1��K��ml�N�EA����tP�!�:�%��Ӝ�ҡ�O�:YZ:���#R���1%��)p�1(A�Gֻd���q�$Gq#�rkv�;�|a`<���0V�d�+�{������o�q��
��T��os���n��>�)p!�#B�:�F|Z��2��U�55ʰ���#/�B��g��W&״.���$��DШ�Z��lS��m�V�*j����g�]h�?$yR�y|�Z���2��g0�4Y>0?Z�TRg��;XpRSyUK��٥VҼ��m�-�"�#���b[L����O��O(�9�쾓�>�^hD�:QGA��KVKv���K��� ��N�,_��3 ���I����z~����r��:�5o��j��Α���\�U�C�#��R�5�NvC��u�����e�B�	����C��r������e@r��nE�Tq(��+"�Qe�*^����t��<lX��*/�'����R�4��ń��4���<�'Z�؋�i�*4M�����_�	*v�lƮ�d#"ǫ�o��#�Ǻ9��:|*J�!"�)���jm��&��9m��e݅;N%>1��)�U���3��i-n
��=i��Oz�p)���|n�!��!����@n`�|�Z����I ������_w:������Or����	|�+C�H~k C �	E��+��w��+��v���+P�����^��A:^)dgYoiD��d+�Pb�����c&�r ��7*-��[��DGu.5X<�)�:��r�;��O�H��Χ]3���&�ϻ�)���
�Dnϩooˤ-��&�o�Ƶ?���+.`��c�c��ȃ%x��C�R�g��-0�p^/l�4�ԕG�vݕ*$c�Y�NW$�EtEz�)��K]Nv���G�7ܞf+x��
F\�-� �
������T�VU
������cȥ�([�Z�f1FBE^^��'l1��ݖjT��J��Q�����Z�N��\�"�ϔ����+�vl��Tq��t9�g�K�G��������$�x�_<\w�wO'D���\�\�<52�����L&���f���s{ȋ3<�|�oR�[ �iQ�H��E��v�<��⦭�>8�P�{y�%���LL5W��n��_�<۪C!�?�¼)����(���lm�3K��^fe�������-��Np���fA�'T�W<0%g'`"�����3x�Q��׫�,�8�ހ��_u�>8ε4,�3钂tT����>�����%�Y���M�5l1* r�������)����C!�P����[�����t'�O�!8����Vi�QJȃ���t�a{X��ǣ�W�O� �ۑ{\�ր�?�d�j����*g���8��/B�=�Q��]�-��3*�d�m��4ä�^xpS�Ns�[�<�C��w�Վ�@���C�؇|�❃W�Ay��&���÷)�c˂�����G 9��m��p9N��:$G��^�W6�4mc�
��pU�2��M5��<���K���>� U��Ѐ�G��b�Ř����(X�����c[O�մ�@@߆G��/�pr�~�3QƯ&�,j�y��s��Z�{�I �S��F�Fċ�Y'IOQG�M�(����",����$�)�!a{���PgU�-��|74�lV	�>�V������e^u|%$�o�R�җߛ�����3q��삿����$��@0�d�ٔ!hC�t'`
᎜����WG3�|�G�ˉ��	}��߾�?N�Aì�
0�)~�0?�+ԁu�E1F�����y�%w�m|�d�܌�37��rq�qJ��k������� �8���6������E��5C�M�_1[K<(<��9����ސ�0S��-���d���G$��waY?~f	V��t����q�-�Yh�H��K��1gO��N7�D����T�c]�VҾ�7��b)QO�����"�ET��L�̂��
V�L"xsӟ�M�_1���^/a'�ߢ�TN����j���p>��1��[/a	Mp2�Ϋ��-��1���N�k��?l&Ҝ�䇙�V���(�v�~�,�Ǔ鉁���[��esBF�����s���eK�<�E��`�C�#��[�I�^��+�kN���A����a�i�-�Ȑ��I(�[љŮ��