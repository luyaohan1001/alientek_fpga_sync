��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1�@�7�bƣ��Õ+|��dδ�R�PM(��~lx�2P��;9�e�b�ʝ��-�3��H�ZҔ|��֑5��؛Q���n�<�M�3�6���&2R��:t�hZ��T�Q�V�)jȫ���ɾ�ZK�|";h����g׵���3�縨�����N'�}?��8!�ګ����=�T�-$�|�J?�[<ʉp9Uϗ`Zp���b��r���H[�<���U�+��?�us�Sg}P��㿖Gqj��>]��H�)�+fϚ�s�j꼏�c�W�ù�M(F��1_��?����q��a3#��� F���b���z��M��E1�`!=��h��L�v�:k�6,�z2��URfgШ�&�̴��AC컨��2�q���*Q���E�����ً/�"�$)���%I�GTҀ��z�X�Ŏ��JC�3}pM��"C������"^dee���M2I̔��/���[�ݻ�#d����峹�i�~�����E�ņg"��ҵ
�F�yu#ӓ�J8+P���'����I2� ]9n����z�3�_t'Q��C`��O�Jh���"K�#�̅H��mvX�v���F�V& Q��=���c��֮tħD��ok�_L0�PD�#�`.���T�7�p��0ծtS��0~�Q���|7�[bA��`�q���VM5�e|ͤ�``���|n��K-������w^�|W��,ǫv��F��h�/32x�*�fQ���O�'Ľ�`�f'�g�v�1���.�N	�7�>Bp�{�`�j��"�������q���[������Ey�7TQ��'F[�8:P�@���a�1�K�2����,�cn?as�8�7���x�W�8�Y��@jX�G��櫞�`�w�:�/�.��9%��Ah�X,�R
�kl[z&�[�$��pO*�j��c�e<���ClӴV��^Y^n���3ȓ����.CΎ^�V1�@N|a��/P<�3�mst�x���?#�����9K������5�IqH=��g_���;�92N���|$'����쓺���^�ŵ��I:�h� �k(�� ŏ���s�j�k&lS'�e�:���Ō�סa��m���TJtZWm�XA���!�
���_�L��3��R���YB_�G��@��:��W�E�/�L�x��
`���FZ,6p=�j~Y��hg��)�o�Hm�^���t�-�� 4$��L����O/���8�+{��9�n(\S'+��h�i}��0Gw`���F��V��*�~���R_~X�`N��Ǜ6B�9`Ε҉��<}}�ۣ�F���<8��⎑<4�3Q��cH3�d�ov� �Sj��D���z(�=���u]�8��ɡ�F�8�E�@�<xjX��ji���ɺG�7u�tF��~cM���J?ֵttCpF5R��E�%1l<��}ZH�Q��U�(y�:A6�G����N�V;>�Vē:��Kg��r[��s}!���M����Zש5�~!V㦓[�'���S����AeP&�)���X�#�KR�ڄ_�l�@���CX�.��LY�b��"k;V~,�����pĺ}O7./��+*w��qD�?5<��f���SlA8���T�
�D2����ë����S��7�摧�<|d�ތ�W�u��\�8->�u)ox<b�c>Z@ЉF��*�k�)�M�+p�r���GZ��5���"?thN���A�^�3?���%�y������>}��T���2IvA�(Dp�� ��F����_/m���a��kt�'�-�d�,����`��g���϶��q�_E)%���d&�<��^�d'�bhi�����Ab}4�>��\�LR�}�����O8���`���fgc�)��ܨv�?b/��4���o�
m�w��PH�0��&S
5!�[�)&o��V�V��m3��zh�������"�Xm��8���m6�P�y[G��1�U>UyX+ZĠ�n>��@�fJ��V�u�O� J׏���/.� �!������W��P��)�K�D-���"���ǿ��ѯ:�<(��)eJ�)c+��XW`>�PS�;t��/0�b�Fz+�c'���B�OM_��Wkdlm
q4�B���,g�2e�v�WC�k���l�M��=��!��f��2�.�I1`�� n8`$��A9���Hp�k���ϳr��3��w32C>�L��$t�O:�܊EП=X�%�F�u�7W�yn�߫����UM�#ԣt��V蒙#]ma���=K'��$Ռ��
��]����.���6M�P�[|������o=�0�_��{��/�5K��R���#Vv^
��gw�4�v���q�����U4um.�%B�"�o�Keh��h�|_��&9�p�V�-��W��0��ɠu�i����(~#P����z �<ƫ��b{9R�_ߕ�w����@�4������ʙ4Dth����@Z�r�!�����Y��@FOQo0qM���%F�Z�I�\L@tVf��~��b��q��"�����
��k������0ɺ�⯂����SKvo�f��)�ם;r� ���k̫-��)��)!G9z����~����ӟ`�IDϛD	�u�x�ۏ�pL��� ��{Ǉ#�!�c?֣�*�.���~��� �{EW��蜜.Ŕ�E���h�ذ�OHD�l&�Wa����k��"�
���8CsU�$%N>�}�1$�X�xEH��Eg�@��W�*���VC�@��yp�lP���֗�[J��t��b!��m�>hkTh�t����6�Dm���dB��c=���N?�����eٺ��Bn���\���؁�6˧/e.�x�^J:�K�Ůo��Փ���e/�Y�L�0����0!�P^[�}מ��8�_�+I��Ё�}�:��~��o��8���JE4��M��H�U�=2�.�2M���U�W@H��$���;�+wr�	��e�gc��G�T0V� 
5����� �B �͑�y��>�)!�QWE��W�lw<��ce��1Mʞ���*z�Ww���ݧ��z�5���&�xe/�Q�UDxE g!�m7��橡fx+c��Ň�Y��t��e�ަ�n$<�9&��	�y����$�!�^��h�}j3f_��?.Hu�
T���rt'&ښ�L����6�w�듇��y7��)�&G�q	������*u��#�*
���w��I7���^&XV5:�6 �(p