��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��������U�5�n�1	�\W��b�1����/�ib�8�GC8(���9'�4[Nw����jO#H�>��WS�JS�_%R�kg=f c�+]l5�����ď2ݳ�s�T���s?�ߑ$1D=kxi�OcT7ϴ�?�T�f�X�k����r���Z	8�Я\�\��y������ơGzb�C;c�?��2��GEPr���4�$E��U_O�>�ѱ��z:X;�%X�{�e��9ۛ_��	�l�y{ba�xq�RܛwD��`T�X�����=6�ER..v[fm?��������^�%��y�X�*H_s���Уf����;:��o�Em�ʺ��q#ұG�G?�o�	t�3��p��=��v���o���M������S��-W���;a��u�-&-�%<�՝7�L�E�_T笊��P��v�B0�ѕY�d �:�H;�#dz��X�~�z��2�p�*�
v����\ &��e��bb}�]���)���D��N��=#�fr{���%::��<�*9����׎Li�3[y��#��*�	�q�㻦���Niв�P�1����T��:gU���R�;��2���LTio��Wbv�ϞAl�K�l1#��a�c~�L4ܶ�$+��g��
X��!����I0I�!��WF��rc�C���؂�º���\��޿Q��b35�����ѵ)d5`�����n��Q����T�[�:����JCg�bB 5��[�uJ�w/�6��!�:u]��]����'ׅ�ߚA	��R��]f�������{$���]�D
]��s���"�b02k�寓���?�8�O���]���GpL�]�����v�q����. ^ۀ�V�����*x�MΏ>A������n��p)��UM��.���=�AE0�J��K>�q�S��WE�Y��R�a� A|����z5 x�
o��:I�[�>��y����
M:��.O���֋P�nh)*X����Coݘ�^@�c���X���Fښ���;T�V��R�Ɛ{y�|�m�w�S<���8&+����H��(W�}MG��p�Lڸa���6
D��b��M�+Y��D9�;"���sg$*��I���T_��-^�����{Z��
���|����Lsw`�B����Y(���C�hޑ�]���q�-����N<��8�<uh0Yj�@OK��Kp3Z�,��y�eV)W�U˫��<�eKW-
��oo���F�Ou+�ߺ��Q�?���a��DT_5�*�v��%1����U�t��Y�,�Bd�~H��F{
r꽷� #]
+�%��i�o�#l,Qb�mV�� �KISN�U����?;+�"^:�DA�1Zf-���+|�?<��9�ۤ��nۏ���s����3k<�&��P:r
d��_
�K��$m}.	�����1?Mo��K��X�WNK�����BC����6�al���3�Q́�*�µ3������� }��s�H����N��"�1�L�������~�����f����PT+�5ު�4��Z������*�X��1wÛ>ь��L�4�p�<E�O����#�C3�I-e�4�u�W�5��g��W6h�T�=ҐQ������4��kU�!�kn`~�J�,I�- ���w�A�.',ljL��S�a��Bu��o�u�����("�W.FL� o�j%'S�t������sW\�̉M�Ca��g_��ҽ�e�ңI� �f�����W �]W�n��p�D��U��V��D'�Ȉ-����%��f�^9w1�Ǉ����j�3��.�r⦏$h��n��d�cB�Ɋ�gl��KpO�!3��t���d���0O���Un۳NV����]k�8fȻ�;�[cC4N�}!^��pI!|6]5b�[�Q��;���E�k�N2�Ldho��t���=��r|�Z�t����6��1�զ}S;���{E{O[���8J ֖Y#�ΰ�/CA��]8�{�b6z�p7OL�)�H��� ǔ���ƞ�k(|w-"�ԗv�������Q�N��
��ٙ\cN6II��p��Q$�a������d	�>0��g0�i�K��	�9��ی�7R.}�ǋ4�3��ހ~&�/%�DvÖP[�̙��v|�a�n�f�[�S�Ad9�N���	�U�<�1�{ɵ��,���$��T(>�����fJLI/ ���E����O� �!C��.{��ۆ�ˁ��K����P�wy[�XQ�u�s�bü1k����1����."��y�$~k��o&n�t��[��A��|0;-��ς�ފ}0N-��
���9�NY�XkW��O|47��I��xC��D�z��4�ޕ^�F� ���F�k��p�u1�Ȯ�)�*?�V��l�h_ΌHU}%�a�"�>t�+Cf��/,�\c�w(?�:?�F-2w޺X7�s(�����h�~�:vj7b���c���|!߂���ءT ��L�d�Y�$��rȇ��y��3��-�}�*� 2��kq�7�����F��s�7����B��)���M��\��g�������9̞X�z�)6\4�����u�6*s��f���刕xe�F��#
gBZO�˯)���6�݄#d�S�mii�} ���se�J_0;d�`A�f�X��7�+�K��B��9��E�7W�,��:Z>Ma����hs�T4�ɇ�A�h#�,6)���r�/��7�{�pj�3x��G�s�ה�7�G�تv��e��?Ե0/�0�
I.G���F\���A�>�#Q6���AfTb]
�r�	Xo�����0�&��P���,x�˦�;^�\�uM����`~�OxD�\/�Ƌ6������A ��*U�z]\x`��MDgg;���w�)�o�ml89��2�,T�p���>!k����Y�UvW|����,��V�P�od�z*��_E/:,H�3]�5��n<�Σ��S9h c3��E���{!t�:�!�P_9��39�Y�9P���1�}�����T��{f�#!4Mq*�҆��-ف��-Xτ����hn
3�f:��X����SGhB7�Ҟ��L�$:�-8%��ҿw�Oi��I�F����ަ�$ۣc�2��6�d���`�dWG���Vg�[ȓ�n�o�%��Mof~º�a�:k���\���}�{�{E��v��u7�&f*���2}�W���9�[�O�҄�����>] *��O`|j-Ú�C�R�J'd����N'Ɇ�-�u�&Ed�;���Ђs��!F8$�|a�y?է� �CK�/��c��6�T�R�9��Nk�A�uz;���;lc�=�E��c�P�;Ae�pUd�[-��_��V��ѝRWڍ}��9�&Ne���QH��G��;Z�)r�j�aD7tF�IO�2�̳�=?��x����Rr�� ������,z�m��R���OU1ה���s�������
J�\"�"���;��m�Km��
��b	�#�s��K�k�>(���n��$,���b�S�\q��+d۞� Z�Ɇ�EQ������
��"v򌵗=�^h�u#`���-�dP|t5����������ȍ$W�)rM������d�����A��e@�]�"�4�k��5qp�O;���	,H��l��x�,���=̆Q�}����#wL�ick��p�������|������0���_�y"c][{Fc0O���y��܁�e��`��\����B�V%�U���U���R)�d��~������|n�a��ޏ xa�F(�f�g�C$X�υ�v�޽
]��S{�.>��)E��\�L�\ᚸ���bH�;��v���O�߳���yx�D�"�p�	�����35���ˌg�I��d�D���8[��8я�gb�w"�0SjL���9�Ү~��0�=s`zx��
���� �1h�9�߮�	��c|m���>�B+'y�?�9�3YyQ��Dh��T��{8aYBIx�G(&6�����w��c����3����� �Y���)��������k�20��w�7�j�N �Q!]�[Lň��尟��Ľ�җ�ꗪ'���b(���Z#;���o�i�nf�VDo�ϳ����H(���
�����Gb& p�7���welZ�t��J>>۶53�5�z�l�E�gZwZ�Y�>���rM�j�	���\z�^�����yn����7���<h�U[}��E/�R�0!�K��Y�>S�λ8������:�%��i�%Qi ��Yb�e�m�����$>+&��v6Z�bY��t�!��r)X���}v� q��'m��=ԘQ�F���S�Dؼl#��~S���0*��O�"9/C���-��8w؄�ȟ'F']����j'}V���ě����Y�[[.gW� s��o�=!m� 7�q�:�?�4&z�����XB?��lQ��*F���F��]O��{���I�R�Y����_�^}<�n=M;�d�ΉBu�E8�>gy:�VUV;����x���%"rj��,�d�y��6c�P̑�� ��A�Y��`$v�Fʁ�E�*0HL��d�A���.��R�c�]�	��z�9�v��n������8r���ճka�	�c�����q�t�Y��L�����
�\-=�/��*wl[@�R��8T��9Q,�7-'���eς]���UE⓼����K�v1`V(���gP��0�zQU�#�!i�o\n�^���qs��k!�>=��ع
���Ɩ�
�X��9��a%���=wv��C3>̖B���ޡ�&J��!����k���\KT���2?܄�?�h���7��������N��I����ٌW+�vB=��|�M���m�O��%g3����ݚ��!��k�-єP���wA{�b���6��� 6�n��BE�3S���K�JC�W�;^D%�\�P\��7݇�K
�8��4+듰��V�9�L�4���o&����� ��"0��S1�d����f������w��|Y��x�%O��,K9_K;�N����aBU0��xd=B^`�,�Oi˲�{��gXʦ�Q+�	1�T�ƕ��KL	���%)�/ �\,�4̿99�l>" �#_X�c��3qϫcu�ш}ˍ��h�9(�_=3z E�"��$D�͢���W-s�F7P���4J"�r�~��jx
���ܞ`�(Ձ�d�-D���{�*O�̸�<�s�vzjOu�H�H�%����؍j0�/�.4�ʹbS��s�Ĭ-��Mq�x��u{�!�/Ek��#Tn!}$���?e��l��,����k�4rەEu����u�Kח+�F5����VG�ߤ;�� �ͪɞ���:4ߺ���u;z^�..?�eWH�xɼ�8�P釈Z	��
HI��w��#+nCrx�W,��Xp�;�]�q �9Tc��M�cN�x$ٯWc~�|@?6ǑcG[pr�D?��%���cԖ��m1J��SFP@cc����+���y|�����<uy�ʲ��#8��&x&�*(�;���ur��m���AOl;G�QJ�<b�,j�+�X:��M��ܐ��hܜ�+v���5�w�\Z�ك2�$�Dm�t�9 u���$�y�8���0͔T�J��M#�y�46�)�89��s2��hm�݋.�ٳ��J����5�3�,�-_���`D�3H���� I|��0û��,Rq�^e�#��L�?�n~��w[W�QTD�̂x>`ܲ:�?�������'������m��e(ߨԎ��~����Z��a+�'�<��v�V�y��a<M �4�z����r<�~�gDU���~^ ���Q,]��:�&+yy{(�]�	B��G랺,�o���v���IǗ¾�~F<)a�^^��x!�	+E�^[�:��:+�]���"�:�^P��Dks�&�Ëd_L�'�a�l݊!98��Z[�-�i�c�[;��}��Cm�%\��оm�����
�o�-�H2c�>,A���a��'�ǒTஎ?�b�������2lr�X��8��44�;�r�UV��x��#�&�Q�C�����s�n���E|.��>�f��b��i��c�;^���!&�/�Rz�E��}$cZH��W]Y��2s��*+�Jī�оM� Z�E�`JB5�^�"Vm*���H%�(��:n����ml�[���Z4�������+%:7���D����F�s<J���R ����+V���p,��ϧ����`���r���\zMp�qa�'߲;4�s�c�3�Q�a�Wyx���䘜J�d�ߎ�%LI䥻�Z��#�\�M��d�G�!�f�����T�0��(��č%���A��5�T;������:P��$��H_��M2.�&�A���鮟�#7��'H�ܴ:H��@�H���V`�:�\�y��3�m7��:nvW��!������a=V���eaf�4V|���J����������H�}�4��rd��S �������|q<���D��b>���]��@�1/����ݥP�q�g=|h��2_w?� ��Q�P\VA*�a�A��%�V`Q
Ⱥ�Ʀ73  qIğ��)}D2\�1rT�d�����m��9��|eR���n�XFG�b~\Y��h�@V�׈��T,���)���߃�3e�$�#�U*&��x� r :�A[zje[�3Ź�q�X�y�3�/�A��~��"��4�6cn���]�Z) ����t�u���;պ��\N�'F���U���ˆ�m3�[����5�U�k�޻*2N�MB�|�;?D���TQ�Ӿ�rئ�$W������6Zo�0ՖW��ѿ54�Z�e�*��ZR���p �>�gJc��+���D�q�4��i��̨����*,�?�>�O1���=B�w�S��GmC�F��
nt��sS`%L.�w� ^����J(m�x�v����G�P1�K�6,���
�м�fj��E
��IӉ��9ej��-o�l-ƉO��bdz��ȅQ%�L��8��w��D����1q|QD�G}�A��	�X�OC֔ۤ/���6��3�k��-{Zx�#0�=��&��wΙ��*P5k[/���E�^{A�2��-6�W&��p\A���&��|��q��������#����]�jh����4�[Ba��#XӒ���H����d���ʣ���u��ڱ�/5whG�5AP����z�u�2*&"�f�Џ��.V� 1q9lk��/|g�
���'$^3̻;��P����H���Q/��
&�Z?�"�5UD���6�~�i 
�cӧ(����S�qʯɸA::��"�;���Y�p����;ys9��F�[�ѹ6��LlEu��mO;�ȗ��r'�ߦ�_(�V��㇃ߠo3c�V�ym��z�#���?�rnO����V���p��}u1�ԭ�|�œ�:�}6� ���>���{�bFH4���Q-�R���p"�³��Ӵ�A��v��[^�#p� �N����P��/pS,��O��Fd`G�'IH	��	J�Je
9���^��X�����F	Q%��*j���Ey��Uk����'���>y�P��4�?_���&y��D��KؤtT(N�?=�$p!q��8��o�J�o-�nY���/��[W��;&y���[���KS�h{���C]�qQ���7G�3c
����}���4���������ZW�����������+�"�\*;9�úE7/�u��4�}O|���Zk��G�f]��	�1��+�2kgk0b�Z�}�`�T��`���5vz��EiMmg��6���JY�T�N��g�9\͎��N��'yޜ֬l�ToF��Ž9�.��q0��,G�]eۙ3��b����-���$C�)=���&�Π(�4�)*w�~���3���9�y"��a�@��[�Z,ǰ�̼7����m��ˊ��A����Xh-C�r��t1(��^� �#�>j��bX�tJ������e\��}u��CI��6W�"<��ld�8%�N�(��l2� �W�bBI�K~���5l�*�����'�}���S���V����+�! c��ٯj�̐bF�4���C���Q~�1�2 ���3��?�g��Q�g�|7��eԗ-�0.��gA���B����qk�%-�WbP�zq�[�/ ������z��b�H�L����9Mj�P1ӡHo2�U̥b��s:Pl�¸�ď�*��~!CMŜ��l�2���C|�ED�T�Q��6aݣ�j��C��ᆤ ��g m顫�X�YTmp�j�b4|r4WOX��)����V���I�7F�����f���c�D����
^��.0d*�Ԋ{���.]�оA� �҈�
�d��<��z�w5Q�����%��t��!"v�����۶嬀�����EP��{ R���=��`
�yGeg�6$��ڍ"Ԅ#�^6	���Gs
Ȳ4�P	�z�1e��+�R�?�}��D�[��)B�M�`+?�����9���l�6�k�Ϯ��RuU<K�H�'8��"F�'���~W��}6�ι�-�p嵘[Oa�w��F���}�A���ݦ1�*��9rm�TY^��)�������Ϻ4(�1C{�۴��9��l��@��w����:�^�٩K���-IG]��rO�?�Qp�p̮�-{����s���A���!�!��Mt(�*jO���r'�A��bD|����?��Ze�6VZ��Z�] ��+�8ux����p~BS��X�Y1{��
#Q�����Wq�S�`�N �� 6���6}<�-����,��SĴpS���B�y���{o�(���T�(�<�Q�~.���k�bh���Y*�~��ģ@sG'���Y�w�˽�3u�@��Vo[�ID�&l/���-+����oc?�XS�b�-�:߸�;)�nH��b�k�x�: �H�n��� )D����`8����ɗl4��ÉnJr���j4�;�8��l0���/��v6��\z47l�s���y�:v���f�ܽ{o��FP�^wĥ"6�X�M�B_�����6��ķps��c1%Bf������k�*G]c�V�w��@iOBU7�u�S�w��1[�?�a��s���9�,���*�fۇ�v,�s�|��n>���S�t��[.�ʂe��ۙ�);��vʈ۷"Q��!>�M�r�V�O����8�%��}o�P���;�v0�#�DlB���E~ؿ��x�v�?�)ɉ����P��+T����=�@����U����SC�7/����}f��8}�O��:k?����M��e=2� 
�M�q�'$�im�"O����$�N}��3�+	�xFj �/9|y~:�	R�s.�����xR։Ǧ?U��ض\�K����BH��Ӿ��͞����۝D%�V�FY��A�zΡCR@�XOua��)J�P_Σ"�T��9��[�G�v���0���rf�=�ߟ�yL�f� _