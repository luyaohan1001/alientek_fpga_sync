//****************************************Copyright (c)***********************************//
//技术支持：www.openedv.com
//淘宝店铺：http://openedv.taobao.com 
//关注微信公众平台微信号："正点原子"，免费获取FPGA & STM32资料。
//版权所有，盗版必究。
//Copyright(C) 正点原子 2018-2028
//All rights reserved	                               
//----------------------------------------------------------------------------------------
// File name:           lcd_driver
// Last modified Date:  2018/11/2 11:12:36
// Last Version:        V1.1
// Descriptions:        RGB LCD驱动
//----------------------------------------------------------------------------------------
// Created by:          正点原子
// Created date:        2018/1/29 10:55:56
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
// Modified by:		    正点原子
// Modified date:	    2018/1/30 11:12:36
// Version:			    V1.1
// Descriptions:	    RGB LCD驱动
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module lcd_disply(
    input              lcd_clk,      //lcd模块驱动时钟
    input              sys_rst_n,    //复位信号
    //RGB LCD接口                             
    input      [ 10:0] pixel_xpos,   //像素点横坐标
    input      [ 10:0] pixel_ypos,   //像素点纵坐标 
    input      [15:0]  ID_lcd ,      //LCD的ID   
    input      [15:0]  rd_data,      //图像像素值
    input      [12:0]  rd_h_pixel,   //摄像头输出的水平方向分辨率 
    output reg [15:0]  pixel_data    //像素点数据,
    ); 

//LCD的ID
parameter  ID_4342 =   0;
parameter  ID_7084 =   1;
parameter  ID_7016 =   2;
parameter  ID_1018 =   5;
parameter  ID_4384 =   4;
//颜色定义
localparam RED    = 16'b11111_000000_00000;     //字符颜色
localparam BLUE   = 16'b00000_000000_11111;     //字符区域背景色
localparam BLACK  = 16'b00000_000000_00000;     //屏幕背景色  
//reg define                                    
reg  [63:0]  char0[15:0];                       //字符数组0
reg  [63:0]  char1[15:0];                       //字符数组1
reg  [127:0] char2[32:0];                       //字符数组2
reg  [127:0] char3[32:0];                       //字符数组3

//给字符数组0的赋值：OV5640 0 (16*64)
always @(posedge lcd_clk) begin
    char0[0]  <= 64'h0000000000000000      ;
    char0[1]  <= 64'h0000000000000000      ;
    char0[2]  <= 64'h0000000000000000      ;
    char0[3]  <= 64'h38E77E1804180008      ;
    char0[4]  <= 64'h444240240C240038      ;
    char0[5]  <= 64'h824240400C420008      ;
    char0[6]  <= 64'h8244404014420008      ;
    char0[7]  <= 64'h8224785C24420008      ;
    char0[8]  <= 64'h8224446224420008      ;
    char0[9]  <= 64'h8228024244420008      ;
    char0[10] <= 64'h822802427F420008      ;
    char0[11] <= 64'h8218424204420008      ;
    char0[12] <= 64'h4410442204240008      ;
    char0[13] <= 64'h3810381C1F18003E      ;
    char0[14] <= 64'h0000000000000000      ;
    char0[15] <= 64'h0000000000000000      ;
end

//给字符数组1的赋值: OV5640 1 (16*64)
always @(posedge lcd_clk) begin
    char1[0]  <= 64'h0000000000000000      ;
    char1[1]  <= 64'h0000000000000000      ;
    char1[2]  <= 64'h0000000000000000      ;
    char1[3]  <= 64'h38E77E180418003C      ;
    char1[4]  <= 64'h444240240C240042      ;
    char1[5]  <= 64'h824240400C420042      ;
    char1[6]  <= 64'h8244404014420042      ;
    char1[7]  <= 64'h8224785C24420002      ;
    char1[8]  <= 64'h8224446224420004      ;
    char1[9]  <= 64'h8228024244420008      ;
    char1[10] <= 64'h822802427F420010      ;    
    char1[11] <= 64'h8218424204420020      ;
    char1[12] <= 64'h4410442204240042      ;
    char1[13] <= 64'h3810381C1F18007E      ;
    char1[14] <= 64'h0000000000000000      ;
    char1[15] <= 64'h0000000000000000      ;
end

//给字符数组2的赋值: OV5640 0 (32*128)
always @(posedge lcd_clk) begin                
    char2[0]  <= 128'h00000000000000000000000000000000;
    char2[1]  <= 128'h00000000000000000000000000000000;
    char2[2]  <= 128'h00000000000000000000000000000000;
    char2[3]  <= 128'h00000000000000000000000000000000;
    char2[4]  <= 128'h00000000000000000000000000000000;
    char2[5]  <= 128'h00000000000000000000000000000000;
    char2[6]  <= 128'h03C07C1E0FFC01E0006003C000000080;
    char2[7]  <= 128'h0C30180C0FFC06180060062000000180;
    char2[8]  <= 128'h1818180810000C1800E00C3000001F80;
    char2[9]  <= 128'h100818081000081800E0181800000180;
    char2[10] <= 128'h300C1808100018000160181800000180;
    char2[11] <= 128'h300C0C10100010000160180800000180;
    char2[12] <= 128'h60040C10100010000260300C00000180;
    char2[13] <= 128'h60060C10100030000460300C00000180;
    char2[14] <= 128'h60060C1013E033E00460300C00000180;
    char2[15] <= 128'h60060C20143036300860300C00000180;
    char2[16] <= 128'h60060620181838180860300C00000180;
    char2[17] <= 128'h60060620100838081060300C00000180;
    char2[18] <= 128'h60060620000C300C3060300C00000180;
    char2[19] <= 128'h60060640000C300C2060300C00000180;
    char2[20] <= 128'h60060340000C300C4060300C00000180;
    char2[21] <= 128'h20060340000C300C7FFC300C00000180;
    char2[22] <= 128'h300C0340300C300C0060180800000180;
    char2[23] <= 128'h300C0380300C180C0060181800000180;
    char2[24] <= 128'h10080180201818080060181800000180;
    char2[25] <= 128'h1818018020180C1800600C3000000180;
    char2[26] <= 128'h0C30010018300E3000600620000003C0;
    char2[27] <= 128'h03C0010007C003E003FC03C000001FF8;
    char2[28] <= 128'h00000000000000000000000000000000;
    char2[29] <= 128'h00000000000000000000000000000000;
    char2[30] <= 128'h00000000000000000000000000000000;
    char2[31] <= 128'h00000000000000000000000000000000;
end

//给字符数组3的赋值: OV5640 1 (32*128)
always @(posedge lcd_clk) begin                
    char3[0]  <= 128'h00000000000000000000000000000000;
    char3[1]  <= 128'h00000000000000000000000000000000;
    char3[2]  <= 128'h00000000000000000000000000000000;
    char3[3]  <= 128'h00000000000000000000000000000000;
    char3[4]  <= 128'h00000000000000000000000000000000;
    char3[5]  <= 128'h00000000000000000000000000000000;
    char3[6]  <= 128'h03C07C1E0FFC01E0006003C0000007E0;
    char3[7]  <= 128'h0C30180C0FFC06180060062000000838;
    char3[8]  <= 128'h1818180810000C1800E00C3000001018;
    char3[9]  <= 128'h100818081000081800E018180000200C;
    char3[10] <= 128'h300C180810001800016018180000200C;
    char3[11] <= 128'h300C0C1010001000016018080000300C;
    char3[12] <= 128'h60040C10100010000260300C0000300C;
    char3[13] <= 128'h60060C10100030000460300C0000000C;
    char3[14] <= 128'h60060C1013E033E00460300C00000018;
    char3[15] <= 128'h60060C20143036300860300C00000018;
    char3[16] <= 128'h60060620181838180860300C00000030;
    char3[17] <= 128'h60060620100838081060300C00000060;
    char3[18] <= 128'h60060620000C300C3060300C000000C0;
    char3[19] <= 128'h60060640000C300C2060300C00000180;
    char3[20] <= 128'h60060340000C300C4060300C00000300;
    char3[21] <= 128'h20060340000C300C7FFC300C00000200;
    char3[22] <= 128'h300C0340300C300C0060180800000404;
    char3[23] <= 128'h300C0380300C180C0060181800000804;
    char3[24] <= 128'h10080180201818080060181800001004;
    char3[25] <= 128'h1818018020180C1800600C300000200C;
    char3[26] <= 128'h0C30010018300E300060062000003FF8;
    char3[27] <= 128'h03C0010007C003E003FC03C000003FF8;
    char3[28] <= 128'h00000000000000000000000000000000;
    char3[29] <= 128'h00000000000000000000000000000000;
    char3[30] <= 128'h00000000000000000000000000000000;
    char3[31] <= 128'h00000000000000000000000000000000;                                 
end

//显示逻辑判断
always@(*) begin
    if(ID_lcd ==ID_4342 && pixel_ypos >= 0 && pixel_ypos < 17 )begin
        if(pixel_xpos >= 88 && pixel_xpos < 152   )begin
            if(char0[pixel_ypos][63-(pixel_xpos - 88)])
                pixel_data =BLUE;
            else
                pixel_data = 0;
        end
        else if(pixel_xpos >= 328 && pixel_xpos < 392 )begin
            if(char1[pixel_ypos][63-(pixel_xpos - 328)])
                pixel_data =BLUE;
            else
                pixel_data = 0;
        end
        else
            pixel_data=0;
    end
    else if (ID_lcd !=ID_4342 && pixel_ypos >= 0 && pixel_ypos < 33)begin
        if(pixel_xpos < (rd_h_pixel[12:2]+64) 
        && pixel_xpos >= (rd_h_pixel[12:2]-64) )begin
            if(char2[pixel_ypos][127-(pixel_xpos-rd_h_pixel[12:2]+64)])
                pixel_data =BLUE;
            else
               pixel_data = rd_data;
        end
        else if(pixel_xpos < (rd_h_pixel[12:2]*3+64)
        && pixel_xpos >= (rd_h_pixel[12:2]*3-64))begin
            if(char3[pixel_ypos][63-pixel_xpos+(rd_h_pixel[12:2])*3])
                pixel_data =BLUE;
            else
                pixel_data = rd_data;
        end
        else
            pixel_data = rd_data;
    end       
    else
        pixel_data = rd_data;
end

endmodule
