��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1eO.�l6�?i~��G!�3���S��u��\B�B��6���g/L��{M�cd1C�q�A��T�O+��1��J�|5v�-�/l]}��/~�kdV��'�8`XX*V�[$Xk)��g�5bLI��m�W�oauc1z"b�b�>Go��#E��I�ϲG0g!( ���Wd��`�a���(0\���̄&M���!;Yu9ĤHfn�g��ݐ�_p�WE��O#	��-�~��J���y����#��_�h���4]���'��(+K��)�h�NKa����Jڥ{���~A,^?ޞ�=:�t��^wO�GA��t���z	��l�����H�o�c\`��r�l������%��t��:�4]�)�A����^/z�e�w[o���ӻ:��	b[���y�ë�ޱ1�R�{�D��8�Du t�iD�{rvv;�t�Ȅ�&���y�ō�?���/���,��#��I�m�H}��������q�Vp�`�����h?[�y��a�H�J����$�!���+��Fk�Z��<̶��r\z�͇R�/�p�\�� L$ �9Gk�L@�]J��d���M�*��q�J��1��1�ɲ=�|0�C%�ߓ-9����W���P��"��@m��*��
E6 �vV?s{�p݀��#*o�nf�g��t�]b̑��A�*!�����.�T雸Q3�JW$.c�ȅ5Y!�����L���2��|�$���Wn�8Tf�B��U�$윋_g d�����sy�M0��3d4���k���]�;Q���.3h�9B<�p_�Ϝ�������Ǣ;�Q�%������w[��g$���i�=������Va_��X�y�GC����r$�Z���z���X2Up1�eĆa�X��AL��`E��$~M���6�N�wR/�]OiH�1_o�[��ڈŦ4�_K�T���҄-�o��H&a�g�i�%<�7�Ql˃I�>�iReN�#�ū?�tzET�(%���zK=?7��9fl�Y��6��>���v$߾va�W�ѓ��k�T<��ɳ��E2�H����)&[P�"���K��g���� k�m�AR`��x��.d
�2'+a�\3{�C���������r���C��<��5���'v���P�y��o�#�b�|)��e���ptD,���!1n
�k��;�F�f�=�&r�3�BN�B�B���Ǎ,�6S`8;NE+n�V����g`�Au=��Ҩ.������E�g#TYoe��@�	̵�HU#��w�ם��(���A�	`Lg�Z��g���,�H ��U�D���3���s����f~1X��w��L_�R̗�#�tk����ISF����,.�e���#y����䈉����e�4�~�H~�º%ǆI�*�Tm?����S��lMRQ�<�RD�zϒB&kx�m%���~s��\;u�����ߍ��dmsUeD��u�c��>��(�x�}��c��M�Ë��?��H����E��K�BZ]���Ϭ_o^@��	� 	O��N|���yS{Z��+�\VkT�*�EU/��f��f��׻����id�$mp"˓�&��^��G U��4�>�$��� ϧzH�	�Qp;��ɣ�
J���t��v��0p+?�J]�ZKk�t%�yw+�^�ru�r�K���1`*_����Af��o7a�����,���t�������W:��W5^��(�#y�'��7R���Ɯ����%I�s�[����w��W+=�G�L�*Q{���4���I70ׯ�{��T��C�.VJLg�\�������N3k�����gZ(�)�O3�Vr��f��@���N�B(05[�1�ޯ�۴��_��nw�QuP��֬���i����L)6`ǲ�h��nؠ��I�ʗ$�.<���Ҹ\g*���@��]�܄:-�'*Һ$��j~�6��T�3�/jY�U\��s�5/y:D��'ZaB+��(��\���E1tK�J��Z�'�@d!*��]���#4��'D"#����^ȫ���妣BH�@�3i+v[�ӫAP���DF��[�Z;Ue]s,���0:�������g`)T%uWg��r΢�����_���Cn�8��h�Ȃj� I�c�F��q( (%�9��,��$/�X@{���O�~j��?�P/q��%�Q�6�[��N� k��Y��R���2�E�}�-!P/�� ���=�*̢e(]�Lvm�|�
��iE�2��;�m=4yǯ���[8�K��-i���	��Ѫ�,��6>�і��޺�gk2��N
\ܙv7u���ʰ�Рn�Mq��I(�ɥ8����A`�J���o6��)ΙH���uǚ��@�-ւq",�fQ��}UG�@��*�����T�H�����;)_�Zj�F5_ª:�[��?�k���L63b��.H�|��`��)"4zK�����oQ�{Q��,g��g�T������z����*���4�����#Ơ�:�M�x�轘x��
���ւ�â~���#�-�pWu���n�'rc�b��h�y��V��mRB��Dgg�SN��-x�K��~SE#�@��.6�����ה_DY�U��T2S��9{�n��i	X{���U�ӊ���7.���e�⛣��,`/YI:R�nrn���x�a�%g������H���/ùc��~CQ������ �,]���<D4��q��6p^HdXJ;P ����7K��)�������COWN2��_,���$�n��P���v%�;(X?�`|����23�m{k��珇��\��z:�[ʢ��<(WP�@��0��棦E�1����#2W88<���5�D3E ��p��`,�(ah[�G��3�����e}��d�sH.MP���T��d�x_9�E��T ���>{,,u�L�t/��@2�>��h��	b�M9A{���0ϵ�f��-�9����0�{s�sK��y�_���R:{�}����4��[ �R�( ݋}��`j���F!fea�Բ�Ea��17��Jx?=(+{UDd96�����VP�x@�o:/���e�k41�����Y3Y?>���Ujߦ4
Eڷ�-tr �DG��R��7j�R��׊���y���/I�|�^��K� ��:��y+Rk����S����
�C�@ ]�	�":�-!�aFB͂�a�?��&ix����+���ؒcÆ��W�w��a_ztw��)�x�"ψ�j6���P�4�E��x^~�������	p-K�xQ�ilsFR;���H���