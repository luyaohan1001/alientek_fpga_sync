��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G�����������b�xo=_�t|�s�o�޾��i:�9�-KO(�I���U���:�K9X	���N[̘�q�R!��H��Z1T�s��DU��:Ӛ��y5 B|� ��W d�{RJ�q��.ie�������[�kt�C��vi�c�0�*��|D����)F�������%�^�|U��v;Ƒa��>уlz\o��������^�bǞˊ�ҡ��UJh�V�D��!��#;=g��|��9��J~����"�����&����aT�?��/#�*E�'��������.! '���5)O�A*�;΍Y�@�Ojҳ.�s��p#�T�*AZ�O���d���ٗR@^L��v0K_扙���JM��C��4�lx�?
�.��f06JqH�ž�yͷ���l�R(g5�x��D	�i�������=U��%�k���RZ�sM@���~�p���g���ڕQyI��6�C�+��K���Zxi��k��;�.�c�.���� |��&W�SO�+��x֥�_l��_!����#�T&���Qt�]H��p��S��S��G�~�}oEX~EYA;����Rj�[̵�o�.���|�7Eh�F��b��9'��k05���)�w��8�$,YOS%�`�D���Ma���}���\b׫DbfPo9�(-��C�]=hF�y���Y)�KP���h ���'3��E��}���؋�y���٩[�9�3����o#϶��Q�F�v��f��c �lM�xT�sP��i��W�"�lUOű?�A���D6��֐?��Z@�
^b�ٗ�aǔ�
������O;��b�"ڀ��69��������$$� ����]<v�(ygPE3!׭�]ˡ僇�):u�E�AX�#wZ���r��������,��R���,��*@��R%��@!Y��ϲ� I�`�eZuZ�q�܍@M_��>��GXЍ�tg�:1�8�����(V�H�������|��&�i��`C{�����(�Y�^T��d���@�5���c�z��ZpGjo>�]m�c�=�0�����0O�n�ac�pfV|D�үƓ<_��ǯ��B[͡�K�~����A����T"#lt9g�8c�o?J:��U1�%�^�<l�����&���Bx2�f�(�,��j �<�'�&)b?�j���|\l���@0�H�K�=�b�� |��l�vQQĞА��N\ ���M���y�ѝ]�`FT�"O�Bn�'�l�ɬXR�`+b�W~��a`���n�p }�U�}QsA�0ĪXP���W�'��MY$�����$�zx�����V����vsaG%�y��\�Lf���w�����̲�!���6�O�ҤN��Zi�A��B����8/�J�d[mh�JC�ߵ㑗hf�ޔ��r���̚z��xQ�

8�ZO-f�5B������Պ=*ͦ6�a����]�3�ȋ��0����J:��;�@���k����U���T�+b�e�&�`�ԯoL�:��ɤ��0��� 8Y��p!�0O�� ���U�7F������F���9�5>ЪS������S)ܐ=���؂��K��u	'����� ��Ԙ��,�����d�J�Bx��W�VD~z�(^4ݭ��;��o�[�Ղ�����O�7�}K��`f��|�F�4�/tY��7�2~��4���/�!ʼ�7��K�~Օ��f)�޼�H��G n��f�h^'U_�1��e�1�p�R.���Km�m�L�X�.U�S��}}�|S�e�s�05{E �ႎ�%�z#������p0��?�Q��pЯA��QqL4�l[�x�f�R��PF���f��2��	,C1�K2 Az�NUq���DS�h�8�~�J�Heȗ��T}w��ҝ�1��ڹG4��s�@�Ӫ�ſт�7aE���8�g 2�����Q-0��np��Q6���2�hx��{wM��X�����5�Nɓ���Z��ą[�����8�٥�jE�x|2'�$��s���I�����~���l<�S�ۄ�I��*�u��+~0�c�h֩Y>��3�ѷ��P��k+�e�$#3Y�F���%�*]���pߪ��}�2��L�K���񝀊#�-�V�-���������N7�rŷ3�Cu�\�kPR�\:�p��˫z�p��!���ʿ�񏜹� u��O-�j�/?S/V}��2����V�U��K|kjn���g+
���N̴�_�5���&�ѿ�פVl�T�������u��ur�7p�;��&8p�� # �+��L#N��֛C����*׍pZ� ~��Xe'�>�U,������Iu��Y1�@����d%���~��(�VPl��Al��������u���Ǘ��v��	;�m��7�Z�:ﳐ���t��e<}��2�0�z���N��<�l_%m+O�c6��h�^�`mё�Q�,�!�Ώ�wqrj�Q��G�V�~�=!!���Q����lvR�������1�C�L�K�5����}=v]�ͣڄ�R������(�6���wU�s:�����F�~�}т�6����^Y�X��z�$��d�o�'dڱ	�1��l��Vv�P-[����0��@��ݼ̀�c�^|7T���ud:�X3m'����H��	̵����W X������N�5h����{ƓKkFCP��U����H��8^��>e#�e��S�51���l����.�^�L��v�{Ӣ�<T��5����}�2.���ְ*�\��f��z��17O��q�����yZ��������P����A��i�`C_�_��
�BE(1dY��f��e�,wM�B�j:�?yu���LMD�ë�$0[H<p4�)b�3�0��=�K����JˆU� r[����*hn�����ˍc��&�h`!,�����#���aJD-�C��n�_4�Z�vH����r1Б��WT���Pc�쟨P9�b�����nڼ&0Z��T/y�.k��z6�4�<�d��$�g4�Gh%3Z�U8�q��Iշ끦�o����wx�`�����c��&�;4�g�ƂT�N��]����f��o,A��o���i�=��"�pvF�
wa�(�]�3!b��
�n�}�f��,uA5-_��M���-���ٲ(���鋬�I�H�w01p*ϛ���%xI���2#:Śm2 i��ދb2���s"��'�%��1�.6�Ǩ;:�6Rx��(�dL�5��NK��	�,��i5�ٽ�c*�R'8��{|�=��X��Z�|]��\4T�lFI����i`�L>���<��,S'����Vr����6����]�Y2��h�C�-�xQ �pb�D�t&��a[
h���7 �fF}��煦��?�DT�7s_P�0c���������*St��E3��-�]&��������UnVm3G��UK����L��W�|�::x�mU�����G3VM�W9*����T�Y�P�/���ݦ�F��Y�����U�,9O%��vel�N��P�L�������ZV�#P\
������C1J7,�Mȼ�X'9��⺢*g�+!�!*��%�	3�+#Oz�P��=�r6�e�6��V��^jf��d5c]p��ګlo��i�+S�+K�>6oC��F� �o K̃�y���e���=�}]�0���)mn[��?����%�ɝ�v�=�$.(�y�E
�/vM�-B������mQ�����:�Č�]���Y�x��P�bg�3R��i�-L�
�FfO2;���K�������|=����zI;��+�����R/i"	g��H!�젠���A<��`$~$��k���8��sC�f�aD�ty'�a�:�e������<l��O�u��!i���5�����&�n�}؉��+Ip�3r��a,���`�>#3�=N b�ׄ=}I�u�Ɍ�#:*�ع��'?f��M>�Paa�g��q�0��v��^�o	�@m�m�Z#�EI�׽��P���F���<"B0���~� �n � �;��?�gO��A�W�D�Jɪ��6� ��Ɩ�*^����Ç~.}�ݾ� ��w7�y�̿��~�xAV��2��b���uJos������A;�P�|�k�S�E�����de]���<+|�|�D�g��+ �䉔��=.�.�T�ɣ�E��L)5V#-�ԮiX)  �IwI8o������1���jK�.W��+Y:�b�`����լp��E�&k�Y�O;�+nj�o0(��� ֒ ���@�n���P���]F���k���;��ʁd.�}ޗ���R9�G�1_g��y6!b��z.�����x������c}�>�{�ϝn��'Ckֶ��ֵ���'�1@�c�jIPt��+���' �g��IM���Xn�Xc*�˰yaﻶӨ
�N =r�[�:�A����Zʪ�r.[_rC�t�ex��>O�T�X�/(������%����K�%U��D�3��J�Ѹ�����ǳ��FH���(V��v�{Ebʷ��E��?Ѣ,C����V�!3�-��K���������LS�|�)���/��f�5���E=�X?e�|`e��+<��J���I���:�fj�(�z�Ԟ���X�7��q�r��~��\,���	���$Ǵ�
��H��/@�|�F"��������
b@݃�yn{�n�����g���U�a��H_��A|P L|Al�ߍ��TnR�ݦ(є�K�NR�R@�
۶�G���r�ʮbE@1�0Ƽ��V雄q��b�c��,7�� W��3e��U"��b�/I`"��'�3���\ۀ�S�:��*s�V[����<f�T�(5o�v�nq��#����
"کQ%�WŔ���������6�+g>�>��Ϋ�oJ�������')�GD�C�N�Tp�^�_)��ɒ/RTm��'�V��n�H����jpe^�ߪ���v� Vݔ���E�K���:��
x+(��R��K���#,������?s��i"6�3e{����`u��M�e�9m,�����又w�z!�t(��#g����E�`0�|�x�N%[�mm��MƼT6ǵV�f;]Ի�
�I���o����ߺ�d<b�g��� "�Xb� �6��E�nW�ެ���ȫ��ߵ�s�w�q(S���^�lV��\�Nb)���\�#zAh��y��4w&�CK�t�t�
��r�%������^g���>e�~�Z��y3[
Я��Φpȩ�8k����մ��߇�@��Z�p�|l`��96ƍ��A}�Pf�2��`�ăUe��1�]��.�%cO���q�+PS�R	>o�n�?�ƽ}-��y��r��&����㭛�D#�؜��O� D����0��
�/瓥�d�\G�^��^Rc�!����'#0Ff8�'��)`J�la�d����t:n�x�km�����H�	��h\
���}�H����9���"�� *-a	�&��.[�ݻ��D2�ꁒ�FD���]�$��ꓱ�4
w�b���%���CB��^���-nq^e���Z����څ���Y��+3
�WTr�,���2�M�F���S^:�XR=	����)�|��#Cj�3�@��|o�}�3��:lo����ϝ��W�
1�qT�����''���� ��RA{!r�%v�P���kI��]X�г� `43��GN�S��<�O�N �F΀#�֩sX���҄�RcAX��O�#}��}j��N���\�|��$�O�,�U��wU�m�[o]���u�I�N'D��v�����ƄsaQ�Z�
Y�s
�SR �Et���æGv��@�W~䇎=�EdR�s��ت��X�k�nH�	]x�)ԗE�/���n鐱&�3�`�o�A ]N�Ռ_r���5xk6��@��z��d,�ޡ�:A��q�<��x�I��+�)����(�����1�����q,�rb���F�q��%�����:�'�Z�KE(�A�vH�!$&~-�b��xɪA���6�N�?}�c�m�)�Ud��}������[�W'���� ~s����,�\
5x����׵�W�(Y��ݗ�u{�Ry�!w����Ȧ1)�,zeR��r凬���W��b�|�@@��:tz�gR�%#q� ��P�ц�������A+Z+�-c,��:ǲ��n�n�,rK����ǿ�z�N�p�F�v�#@n9Q5�eQ��hm��iׁ�7Z�o�ʺ��oK��{���-1�ph�F�%N�x�l#%κ��|��a����|���r��=rH"�1� ���5#iEI&|�dZ6*JXI,J�-C䨼ݩa8�"4��_	�c>�%}�U�d���姶]�R2����x���AHs0~�e�E�v�:�9f�^S�/K������PHS�U"?:W�ڴ��έQ�A0��2���K��-j����Oo�1s5���� �"�W_�5�S�Y6Qw� �x������WD�� ��G��&:rr�W`��d�߭*i���SLg��*�EGq���XsoW~T�U<�D$�?�+��yW3i�ev��m_�
e��*h��Hl�����՞�l�6� �<e���$q�E��#�4����xI4����c��Fo���I��S�e�ν�3�;��e��L�k��C���5��-��b��Vq���Yc�vӤ��$���X��7v[Q��Y�:��s����#�G��m�^�X�![W���&����hGA�ޝ&b�8O(u��M|gd��'8l�rS���?�}�do#�!GD*�g�	��ad��S���͒���9��JD�\�0C7A��qWIч>
/�ו��(����,��͔�O9�����X���zj�eK���2��@�r�:��Io(�T��x�����lc�kẽ?�T��a4I�T�9�S*I=_2��v-�$����� ��y�m�Fo��ߝ�;�hLy�|��>�!��i��(MUA]�e�p�(�K��Ƚ�}�g��]r[A����}Lap!���Qԗ3�h�2�4%>V�j�I��=����ɅHe���\���`sR��M�=�:�l.��N0���)w����̾�|��ڼ�Hr^huf��^���eo���	M_��8��۷�<A9�eU�Q�\�nb��2W"g
�k-���P�c�>�[C>m��;���)�:�s:��[�?�˱��Jp�E�r�����^��b��L�%E��c�$�6�TTPh;�t��p@+텢�;1�o�w�q��
A���##O���V�sl�m���I�]� �y�d�w�?~��G5�yǛ��86�g�K{-�.�:r���|�Uh��3�<�h�(^ʛ����=�7�F�=Q�ޮ���L��N̉o�Mh��K'�!��,�q$,Ok��[Uvd(u�R�̖�Ef�ݎ���i�cjM�0SR�Jo��3R���!, _�m(��4O�ր�+�I��Y�,6$Y��>�I�9=���\S
���vS���r�@Ā�����O*ϣ梹 �N��<�cڀc�s�[UMgvzq��@��_���ȴ@�iOr
���	^;����ވ���*���=ͷA@:&�x|�:�;�C߇�9'g|*�]��)��Fy�?�;��i��kj����.&@[�Zbwyύq%{�c�H��dr�2��d0\XA��tTy�1���Ž��m)�� �"k6�g�htE")���߭�sH(�y�/����[D��8��R�.W���9hv�dŭ�?��W\D��(���6>\U?�ZPA�C���I�P�_�ظ6�.c���.��,*}�s�i�:����J1��Yj��Pl�* <��I�FN��b���
M�3P�\���4-���<�&E�e3h{H[
ߍ'Pe@�VX� r_��d���f{��}��;��*�:�σ[��׫ޯ"�����I��O��kqR	\Aɉm�s1DOI�%�Lf�WZ̆rg��^)�s��NwI���E��>��S+��	_P >8bW�����?��W{l��A�D5��_i^��-�X��*$;j0��>v� I�`1qu"��k>��O�$4�X���&��v���Zw���)w�^����G�M8���r��(uu�I}���hʛ�c�Xc�SN(��rw��ѕ!��f� ��U3��©?�c�/ʄq*>$���6?�/��'�s�࠽Cϼ�����K�� ʊnޘ�~B�]�����6=��1�J;��#�4(����7��0/��#g�p`���V��o�]���hQ���C��>kT����m�j��;��{<DCL�A@��G�O
��J�E>�n��Vm(��
�i�0�M02R�`�+�{�F�Z_
!�o��&�%*F��3����	��x�;��ojv�I�~Nt����b��܊$�xV��,�	��T�2�	�,a��
 '���>���|���܎˲�BF!I~��؞6CE���#�^�vL�-z�̝�qa+�]�yE�K?ԣ�qP8S)U��?)�2�Z��i+��]�%��L�Ɏ)�����!�G�/rIo6̫��@ϸ���|���4:������[B�ޏ�sw)rTtV=�Ik�T� 7�nI��G�K@C,�)����1?ia��o�0�*�8������"�IV�5��WXh�N5ɾp�?>�i�NiaӁ��
��|�Ҟ"Cy#��r�x�
l��^ 
p@�_Hy_H�3圗��Vn��"�;����C\���bR��f�Q'c@�2�M���t���ᩏ��K���/ ���T�s�$��7�U]�1V{x&����sOG��=B���4�u5�,P���b�#��gs��;�ߢǋ��*�G��4ɝ����vcR�쩡����O��ǅ���X���"t�kK8�T��C�F�kJ*�N#V݄g�F1F�s��i���W;?��ؑ4�4�>�^m-�_�����ܺ#��z��Q�Vy@�RU�X�$Z��������)2��z)�U����4H�����oW��F�H����/������*�v�\����+@�_�Hv��¤�~�5�,[�2�O�]u�)^���g��}9D�ɐ
r��/=���-,�� @l+��K�Be��Į�ջ-h۱����0�ޝK�T����	`?�I�-�R �L�b�Tp4W���!Y#P�ݬ�����d���R�V�j6�Ag��2)��,��]�y��IrUd0U�q��=X�L^�He3��<=
v�_���)8����S��`��>�g��˲�����&j6^#Dy;�YgR�����z�`���eM�Kn툷6cF$�BLz���U]h�0o������t� �W���Ø���t�k�C��������8u�^��B|x�T��ιS�����Ov��7.�+0���(��֞5�G0N��H�҈}�Q�;^5n�4{1����x�])��O0�� O�E,A=j�����k��w��#��8�C�R�v8p�*tPD�4�2v�Yv��%���<�b��l
�Jo�������e�u1��k=�A{�>W(��	ffأ����@^0����J[���`�q�9�!���
�	���h=��7R��Y=E�c�%���n��P������SJ9z���%���+�E%���=�@#���*ݽ3O#�2��Ѿ�$wU���t�g<��`?��
{�`���չ�GخU'�z�(y
�gI(�I� �-��'�JQ0�Ka�&h����=�v�W����H^����`e��X�P�J����{pR�'> K�1:��`���{˿��:&n+L��qsH��Z����0AH��;�,�A��3 k�R��������z�� �A,:@!���>�Nʡ':���Tû���Ц����g�Dٹ��B�1��}��E��v,�OD� �Y�N��4sb%]f�`˓��� ��?����?�ys��h!>c� �G�UD�_��ϭ��;:��\�^�\�?�~-j�t6�
�\R*|����G��`I��t�+�3��wec��w�'�CM{ob����Фrs��1'wù-�k�,���ܾ9灬B�*v44��e�!�v��I�R���(�|�.slOeu|�i�ғ��K�P��P��nI&�:���=٦�� M��M�%���6��!ZO�?'�(Ө��2jO]�hj��ڝ.�w��rv8�گNq�;fr9�E�VAP^�m�b*�TbO�v��4iA��@1��?�j�B���i�{�;��K���qx�_�U�8�K���RPss�����͚z�X�pB�LQYz�`��N,���:uV�l=u�jc�3";k#�����ܜ+$��Ƈ�`ւ��I�����ȧ�{k��*Z�m��%,�����ƍk��f�1���Ɲ�溂N+��>)С�[��.!�E^	4����DrR��wo���O�%��t�����n��r�u�,���@���%���qw-wķ�(�E6U����؟���-p(��G�rI���Oa� >��;�ʍ`��g;�I��)6�D�����F3y��yF���6|��M�ؽ)V�Yӿ����>�ƿ0۫#a<��/���o̰�1���a�d�4#�f�\LK���ﱞv��k��0�;7J@�wQw�u*���X�=�0�����ڹ4]�q�k���r����1v��?.�G����CYh�M��ϸ�����Te邨�`�*8=����ּ�&;�NTf��7
�r�n��d�@�F��(�Fˇ���*�]3W :����PW!�"T=�!߭�9��l�w��{��34zH8�k�HY��ڌr�8��$S�ŔM��J(qɎ��xw���)�pu4���`�"�����1���7OX���=�/��p@��`5o��<h�}��)#@b�h4p��V��zIy���(9�#�G��9���*��Y���_@ey�u�Pz>=���։8s�6<����v���-���k�P�� �GEi�( ��c�y��g�h\cit�eی6��\�Yl�\V?~v��S���\W��]|���"��%m��c��H[���"��|�'�
�Zi��C��L�t���2�c�(e��C'	O��ݬ]�9
=���Ge����P�������r����Xy�9~�8&si��;�@r�*��FH\������,<jY"��S8�K�:Q82�_W��Y�5�C���% i>Iq�M�*,�q���a ��
�X� �#5��V� �+�rQ�EU+����[�K�;���;ڀ���Z�̊����L�~GЊ�p�BW��8RJA2���S���k��U#�*%��6}ۼ�̀F�&�/�<��`k�	[��k{�|H
�Hb�P{G����<�b%aF����;�?R�!���j�jY1Q��c�ZNJr �Wc���A6?6��:�Z�b���/�6A)}l���T��!=�%\��5�aл�;ط�][����j.dZ�l]��Cf����z�	1"7���u��t71��w9D�	N&9��H�k�>)������n,��L�����8��Ѹ�|n�/�1Y��$���0�>�S�F��I�]t�h��v�ʕuR�@l;Sg�{+'���ć��ok�6���n��a������TPdL5"�;F��<���Fy�W�|�tN�H�h��5�4����$�����e�>���K�3��χ!xM'�Pfi#km3�I?���K�(K��Ik2(��D�1%�v�6vA䶿O�����m���j�S�n�8�Gz�-�i�V0������jƟ}i0_���y���?�P�#0��TA�]�|DH2�R��h%2� ��x#U�Z����#�4jWX��G�Z[�"^�_䢏m�Ͳ�Ѕ�Z�|b�����ݢ�~X��@dߍ�^R�վps��F�ǐhL��rΥ�M�z<�u��"X���R����.tk�3�� VE>�6밁"��Ts�<�sTHB�Kn�ZdXχ�p���
��L��.Ӊ@�*��H����S<�g������c��m�AQ�k
UYY#��1��v�+:�wa�6�8���V��C��OU��ӇG����>��K�(��5�H�/}��^��)S܁c���`)�8j���gp�)^��d��a�"R 0�B��8 ��5?izp��ze��و��۲��p�q"���kJ"\g�3ZU��	"���7.k?���g�Bە[%pr��V��Sh���_ߴv�>�P�_���Lh�.��R�:�5?��̳慾�>@O��8�8�Mz�����ZV�Q��T��d�`m�^�^1���2��5_��.|u�JL	|O-�_j%:��7���D,��t�6�!������K���"��:�/�P򅶄;����	W�P�1���� ���	|Γ��L�fE�332w<e*GFF��$�v�N�</�yݷ��$�Kۢ` Iw�����������:�k�L�i�������p���`ݟ�9QL����_r�!w$�6˛h��k8"�e��;����|���s�M��)g��=������S�(�H��U��X�wLA��0�T����O@�'B��5�����r�ҹ�ɷ!�g�-���˝�ɠ��	q��y���/���mtq"��iK��s�9k�w|C�س���7i���IbT��[\u��	� ��V�sJJR���s8�չV�����/O̙7^ǀ���q.���y��GA�rn�UZ��%�N:+c^�LCSqpE� ?���(���7����4-��d�ͣ��F����K��3�M��y�dS��H�[iH�T��H�H���'Ah@���K_���BT�W����!�?��W�`8�	uZ\/mn�_�uh|s�7�y�r��!����\���>�(�E�Q�+xm|���A#�ϋ��*��Ô��A����H/�W���aܡ}��l�a2��a>f�>� ����W�h��%_����0�ӡ~1�J��~�����������=`����_�a׃��B2}�Ag ��D�J��{_Dk�"��_��绚�w �k��:g$�~�ʣ0r�f>�Z�7h�K8��*oXU!�_�qg8X�[��{!��/��Ao���uC>q��7�$-�Y�4ݘ��^���Q�~;�q$���K���bz���m�3
ń_yE�c�j6���A�=]^k�BC�̴�1��o|QS��|�����\�q��Y��3o��h�B�?oa?�� �����>{0��uC��9\v��W�wH�x�CV��I����GZ)�A���G���;��N*�3wz.*�Ø'�	�8e\Z0�
;���F\��k���:J�J�x�,NZu�g�F5/e/(1m�G�9�+P~3��S2�;(�/"p{㚨��ԜwK���U}��YUn��kb�̙q�}��[�ƛ���zҷ0���ti���[����`Dz����.�i�&.�ߜ�b��7b�O��d��i�5�����A�$��A�'�s�\�^mg���J�U�T��)� v�p���L?����o��и�6�w6�����+��. �Y�G�)���1k+�k6�蓕@��:��ȁs=��嘺,� �k�<63�ޗX ��kr
L]�"`ś]���Y�5[�o� �0��-�OR��\�~�b���7e�����}E���_�L���E�Q~�V�*�l�B�eQ����̓D	K�������h������II	��M~}$����*28�`
��A@+;]��d*Y|ov��ҙ�g[@3A��R�{�lX<��E����ڑ�������?��g?ZjaZ�#X^u���I;n ���=!I`b�m�b���`iL��[��e���i�YA&�<F�*���M{i��&Pe�˸����$>C)봧T�O�L�=��.����Au����s1�����'��V�	�jguV�O�6��}�ޟ��zB=M�gi5�8�h��x�XgK_N�/�GK�3Dh.�x���n�$|D[ ����Y$��{��
�j� ?���0�w�I���`5��SmA�X��o
��	����D8�a�-�Ape��|re�����8����k���Ĭص*�5���HRϨO�&b�Xs��c8�����N\qX�T�0䂨\M�}A?��ɥk�I8.�b�o��!���E~��n��)|��U��r
@��.�R�G�Ov��z��Oo�Q��*�g5d:�"����Q���X�=�7x�<YZ\��|�c���p��6F0�a�i�`�8��Os>����L�������QM�����A&��b�]�9����%$�!��� �)��UrI4�j�oBE��ԉ�8���:C�Zѳ���������òa>�X�����Hր�Ʊ�OA|����{A�o�_�}/�v\�a8෍�J�#nD�5EI��L��䖚��(�S�m�~�$��8�&MQ���Գt>:��}P��\�֭ɘ�(NKB���q
(diq��$�xW*iE���5���>6�q�eZ	8w���2vz�\Ƭ (@P��3􁡱^5�74���5��������&y��0�7:|Q�eT�oe���C�d'_�,�*	CL%i2ru/F҆��[��[v�"�'��vW�Pͪn/}�8�Z���ν�F}u�	���e���`����ʄp^��Żtae���k�u:���yL�����}3J����_�L��U��`CI�|�ZS��e���K��H���w�*n���`lb��t���	pt�B���ȓ����O��J�D��e'Y?���\���y�?������p�r9�Q�_i�x��IG��qV�ً e��k���2����{��]��%eah?Z�s���/K�.�{
!����/:�ZT��e��7���"���p�J����Q{�5/:��3�o?���!A�1�-	�
�fpC$����[ӏ�F6Lв�r���ܽo=H�*)���%oյ9]2�|<[nt�����Iޱo�(Sxq�H�T�UyE������5�O��=�2$��'� �.o��o�i��>�u;#ӡ��R{�6����p�O$n�^cW��_��S��(�����D��z䙈k+)ϹDٽ�����`���~���g/��&FL��Zip��3ӼS�03V�&���ˑ@6�ũL;D6�mh���<F���	�*�xb�4�N���@�vd���ȀT���!��