��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1YS,�>8�����z9c
�7�\cݰ�g�U��p�뛱Y������%�ü�`��$��p<T����! ,oS<�S��M
T�� u���%���9����+" C��˜���xm�?�����-��WZ��jZަ����D�D9x��yao8'�M���RMԛJO�`��䆄@���#9j.2 ;���c�.P+�lT)���]ִ��2�zo^��Y'�l���(z2�Em�����[RJ\l�� ����Ԇe�5j��mZ�����A7%�� ����Z�./TbN�����w����j�W�(����)��k]f6)��`�j�����j�#Ϟ��~3k��.����֨)`)���&1&��s;(�Ar��H�ԅ��{y>�K�?�zŰ��l�s"a5�L��h�*��R��f��$�5��Cw8(�����D�;��p��m�켷�p-��v��0�cO=��+2+��C�D�Ǎ��v=�K"'Kg�hZ����s,˨dVIX"s\������1��F���"��=��Ra�7I��r@Eى�h�}&�)J��Xm�P�|����6�qC���^�޵����9��Vh�����|6���&Ch_�G�l�S������q�g0M�3����g*�Ϭ� D�}-�$�����{�n]$p�����9�P����}�uEV�%�	�i��0�#��eC_�ǲD�DT,�;m����۝	��5��߯��STK%�� w�6�P�]Ml%m�P_]�������[4�A������dP���`�k�?�dD(FR��68�n�:c$�)P��;b�*�
_%I�ѵ���F�j�OFo�[D���1j�"Y:���T4�G�HN̢z)����^Y/g�Gʠ��]���&Er�w� .�%l'b��B �s��V*X���s?�� �2�7�\�t/ٹ���;�5Oe�ʥM���Z���n^u0�ώ�#l�#�vc�N�$Z+T�������{rco�0C��k����F���J�n�!{�g��F (�_�������ճ@I�
�������F�}�/u� ±��x��p�T��PP�e���pBt�nϔ/�Ҁq��J��-��Y�'��эM 2^"Ҥ��r����hVt����v���.�Z��w�&�b&����ڑ1:��/%���]]���1��=ɼ�݉ �J_�c�!����b:}�|R�ԉ��P����Rw����AQ���jP������`�kF+Gz�t`�j�8�U!mQCMo5��(��w˧�G��&^4cY��,�Y�@����+�. ��z>b#A0'�DH�F1y��A�)Y:Հ��~o���A���1u��!�a�빩��(\}�R�F�E�%nԛCe�&*��C"�*�Y�f<\"*�`���_��g;�~�\��Ƕ'-Le�\Ի�>2&��`X���ԬrR3�|��ݻH��X�R�iU��g���}���u��2�^ƭ6s^-VA�H�k���^
h��K��o+��5z啼��&>`�S��#���r��`�H�v�����D��h�8Z��i�@E���£K_�'~�>O��:���$d�3XMQa�p�[��C���C
Ƕ����Q�R�[�e��4��K`R>�*¨����0��_�(� .~��iW̛"��Ā(Gl&g��U}3ЙA�/Dh�!��P��C�c��Ϙ�?2*�����C'I��'�Rf/ԓ�T��)�K`�R��������&2)��贜�#�ɗ�e���O�� =+���[��Ǩ��BKU(3}췒YX{v�	�_�2SA])`*Oc&U|��y���b�w��Oy� ��}�~�奈�Z�ϫHM^��7�IɘI����cAVН]��`�s�������n��<Mx-)x�ߑ?A��n�}��Mh���=���&�NPh��U�E��'dȍ��ԟ���˴��ji�����/�q�8V�Nm��`B�;ڛ�ۊ*~n��T�����5CaR�{Y�[S���F��00�S)b7/ƪ���^�1Z�����Q�4$��A��9c��s��k������ߒ��T!�Y^�E�2�"V�vJ~�t|��}ĕD#�ҷ3,��by}��:"%��"#%�x�զ�C}��KQI��hU)��"0���6t䏚�/�B��N�_�7neپ���p\�@�]������6~�/�g_B�2�<
=������q@6n0����;���=��]�b	��:���0��BԸcD�!oM�ѫo߿g*�^�kW7I�c�p;ꦒ�9t��ߘU򴗏f@����vP~\8f1������1'C<.�ӡ���#c���h��:y�+&�1��G�o5������ٗ݈�^]VY׈����JŐ`ħ֝i��.�'��c����BA�v:����]�/+,�rHo�m��[Rp�༒�}՗�'aB4YHw#��lv�C���P-եK��
h:�$6�{,��i���J8(�mnF�Ϳ��V� ������F���8��6�D!2�D	���Fb�M�ָZ�m��ȩ>]{F�m��>�G��0�ִ����1�͟���c%.)e�ϙ[����?�]o�9��2s�B�v�ح��kc��2/f�?ZϮ��9!�-?�;��'�>�NWv�/l��˦�=��mgW8Ǭ���ڛb'W�a��$�n�T�({-gV����M��'��m�A��"��ec�
��
\bF�.#��q�).Z��Ӌ�_�m�wI�|����S����"�������&(%NxbY��F|�L��5q���.�k�}��R�:}�>���9Ř����"|l*;t�e�i� W@�u'8�����b�u�3w��E�TS��c�$oZ��--��rպ�E8���A�|
�Tm@l@��}��y[�^��w�� I��#:�>#cm�cE BeD����9���\/�؟M�����J��(����S� '� �P����[���&��2��-���T/�$E�7��������<��kr��wMEhq.�;B�9"�^~	�ڷd���r��\�K����ME���}7st?�Q�����vx,*V�&o�\0O�^�!��.Z��*���H�2�5�[�Pz����u�|5�?~8	�sە�<�U��'$�t��R��C�'x�w;�2��h,A�u:��`U%��I��5�7�67�!�_N��;:ƌˏ<���p!>�FW���[=��E��'7�t��K L����}�3�j���������)�N.ѱ�,�h~2������vp�k�L9<�i��mF�\v�c
%��_(��/8g�7Ǣ&,l��p���ۺw�4���5L-��>��q��_h"�C4J�p)���o�'HaF �Wh��j��[6�z���Zu��V�̈́і��u�uVwjW�/�ثJ��Kmx�V�]hr�k9�ڦ@�x��˗TV�k��ٙ���\h�,��''��^-���g���ܴ����v��k�����l~gE�wK��ޓNA2���/"W滎4�F���o�X�����߼Z�`*X��~��rZ�G
1�/�l�jA��ELv��G�k�F�ߣz�|��]���#_��4r�|�/�s��DQ��C��*tN3�s��9���/@pq���hOcrh���N"^�,l�7EZh9�9��K�v����RC�C'���(�1LGݎu�6�lUA@�������TI>eL���~�@x���k���\�/���i�_3J]����<ႿrqMDZ4����a���Ti��hg������]�^�j@�55�U��Y���#��gj葪�!�T�� A-� �g1��q2s���yq�Y�_lFѮ�L#�f���ݮ"�3��H�M��r�;	Vl���?u[MG��w������f��4�j��kK��wo^]��Ylz�D5@C��K�iI�������l�B(y@�V�+�?K���h�d�:�\����(}�M���۲�˾V��|�8�kR����=I�x���bW��Ғ�RA~b��
�tD�������>�����0����v�)1No����0�Ň���a�&�n�c�&f䊳��>eV�����X�Tg���4�s)�,�~�C���х�v ^z�;����5�\l�Ş�/�e�L�F��_�]%>�D����q;� ;/*[�n����9>����SsoX[�(�Q��l���XeaOT���C�F��2+zE��ng��X!������hI}s������A����q���@�<İ�o����_-���L`V�W�,E)�bp�v<�b�t&I�M��YK`�q��@!m�0:�M�7�'��_�\���6'qF'%y�r�V��Ю2�)��m��ql����.�]���R힬�@�{��_�y�P�g��ڮ���˒#R��i��I��>�7X��&w#�ks!�$ޑ��P�4d8��o[f.B���ObgxX
ȅ�ة�ZY�������:f���&9������s���9�����Y���n�Ak�y���YF\��D��Ǟ�~�C&�[�g�o淀���R����XMȃR4�-O����@�:�}�qX���ď����o��p'lŷ�L��ݒ��8�ڠb�p�1�J���o]v��eg�{�U �>���9��������K�S���}Ě|���+�t�[� �v�2�v:��%�)Gyy1�9���=9lm�ʀ�o[�騇߮��2f�<"��%��6����Y�E+�+G��3��z��@��~���'{+��@fR�G�p���g*�Fz1']�;�j��'�}$��;
�8,�/�����@���/C5���7�r ,zr��Q��&�Ů1�;17���h�f'����sЏ:�gq	�=���笏#�wgf�Y����\X�Й[�FY�\IY����@�<D�ƞ�8^�Q�l��Vg!�G���zL�7䜴;W�\}j�`Roc+DŉtX��m��h��}���x������1e�g�鮞��@'YC��˕	��aS.Ӂ!���L�Qa#��<0H���+���'�L>����Ϙ#dR�S1�����]cx��0�=�'c���sV�Y��vB8[�X�5Z��^Q% 	r&��p�B9��Kjښ��_�5V��8�������3�M��c��W��S�h2e�	��ti�Kd?���Ψ�qrud�@�輖E�2*P
��G{\jC���z���%�y����i�Ib�S��i��[d>����+g��	N�W�z��扽F�%�oI(S�\�	_�&�#�۵�0����y�� �8��87䊥d#��B_>A��JP8���@;����r�Gѕ���6�(�%�7�x^�dX��Ҿ�[r�z|pDU�}����.eN�qGp���%-d�Gnz����[�@�g�����Al=k��ΰ%�V�lv��2�JI��6CS~�h��������btN���xPAeL\�y��~V;"�%E���v�n8"׿�1G�+��O�&4��M�MSEُ�k��Wٳ� Be��X�U�(�����~�*؃��O}� �Gf@%�쯝z�Rs"2����	��`X��aN6G)xB�>���R�A�)AM"�G��A!�����H��e'6"TXԚ)]��OS�%D��3^.;�t�a��l�ҀQ�e��:�U����׍�}����׏8.Yl�������wI�]��[	Zcz~����c]fps��6(Ȃ��f1$٥�������~7̀�:��eA@��	T^��d.�M��Z<O'oDЋ�榶���ѡ�Q^`���C���hF���9F���˘D��Y��Ă��%ϝ3����C�*�\�"��6WTcgS�ga-�cд>�ڣ�?����k�X�S�[	���e�AO:��r���<�F��{�w�V���J}�V�{�S5�v|y����uf�I�)!��-�n<)������o��SNBF��\�S7V��t!�d;E���u����[��í��X�J%!����|����33�`O�z@� ;��S�o󛟐�fԷvd��c/�5�Nڟ�A7�v����"�e=��0b+#)hm���Q�HY��8��4��#>�����P��OK���1 s���85.�ݙ"�T�Wd,+hd�`$]?�9b)���S�5RqaaMp�CaM� =�U�V�G�ŀX1�}��q�(s+:PLl�	�
��R��XF(@ \�-�ejgj�{;#�i�Ƒ�JP�z�s)'��H�o���t�HY���� wb�� v�O��J�E���sne)��1��<з�Pa�9ixB�E�Jv�ա)�H��R�;&	w�����g#kO�*A��O���qHKY��Ҏ��ປ��w����� Y��D�ٷ�ʳt �b��n����rm2��CXۇ�O5[%s��	��(ǈ�`���J5K�DԷ�8h�w��|q�^��E�չ�֩��|X��	��)*��"��\���OZ@{�0f07��(��A]��!��ث��6�$(`	���(������2T�'I����
�����<8�HR�y�x����\��2y-��K;�����f���l��7�g](�C���y�gW�e�[4��&D�Hɬ�/�Fj"�:&�l1߳L9�vyϱ�°��H�2��^�{ƚ4*�,��1�;@˻:_XU�Iз�W����~T꥜3@�e�˩.J��A�(���0�����?sE����+�|H����`�CM�w.p�/�i�2�eG>R��8���?z�G�l��6	`ܷ[�&��W~C�]Vx������b�|�ԯ�2��m�"����] �{����Bn�c7�0�=0M�C�#�Ⱥ�JÐV�kR}0U�~R��g$�'�a`���[k'�&�0�S��F�d�R2`4���ĭ�]�g<��~ȗ��,��-��\�a��wt�	�P�_h2��u���汼�K�WYD��Ӽ��K�TRiä�K߼��*-zj�09�֦	LHFko��Y�8W�@��5҂m�\��B�M��	r���7�܆ϓZ�V�<It}���O��}t�9+8x9�Z�T�!-���1-�/��f(Sp�S���q<C��P/Q�������uK���4�?�dc�l`���� �����fJ�6��P1 Ā�$4�M��pY޲LF���u�QP@[���N�}��H������7'o��{���$�M��v,v[֋l�G{���_y�;[�E�����"���%$;ɼt]	p�:� �ZHd���޹?z*'��	�M)C����~).�ь�����J$k�����o��p�߼w��y��6�M��!q�����+(�L���ʨ$�Yk�����f�ʅ��tғ���0����'l�K�`���5�d�D!r�
�G�a�N��RW7wM�k8��jr�$�������'J���C�u�ُ|L���ѩ�x�Dؖ�|�Mz��@����n��#.�/;1"+2�.������,�s��E{fD��GWuŶ�`~�WqMnֹ�*�ۄ�l��P���o��,�y|��5[�/������0�����Ev�e��A�
����iFwژ����-,AT���hi ZaV��m���y��B�$O?���SH���}f��q� *QX��e�7�f3���Et�Cť�y$P
�G�k�6��:�����;��bl;lHy䨴]*/:b����Yb���2@���C�R�j.Rd_�OJ�ziT���g��AH����ط�m�f���{���?��Z����]J��KBO$v�>�l���?�#⬠z�n��՛���Ej����q�U�,�:������"þ䠞����Or@#�1S�v��)�FX.�L�׊sa���Ҹb��/+l�5𨉳��Y]��!i�U3��sw�����.�Rb�$ �Φd�C�c*���E�M�p��d�Վ"f���H�jĴ�:煾��L�i�*xJ�p�.����7�Ď�<���Ql.4��o�%�n��"�C..)צ
#n�E���EZC��'���5m÷~5-�|7B�����t��q�XH 1�*�ؾ�Z*�sC��T�O�mk ���dD�w���(ݍ��ٍģy?K�b���"�S�" �n�w�^����2m�W
W@T��l�ʣ!򐩜S�#�u(����3&F[�[��"+�����Ѥ`�ER3����=�qs�
⹆��%s����n�-�ޠ�1�x0�"Ȣ#ʌ��bh�|n$�"?�2��ցp��U���kD����I���^��9Evor`u��31@�kcMU�cK�! ߓ 4�!&�9	�,A3͞_jc}�fSF�Vn�gX~���w�`�,�ټ���õ"c[���z��N�b+��������(��b��Z@R�3��!<0CQ/Ƣ�oIՇ��.��Xߥ����!�����jr눗�5{�t��S�p�+I���:*c TI��?���B]���j�O�����N��ՕRm����&?XN�)��q6�7��4�o�X��y���}��������u�|�����W��u��̧�RWB�zji�'�}�!����!I�'�,�͹�;��z!-���g�"N"��J�U�1�6W�b&�.��Izn�^����'�,z�H]�� Jb�l���qbw��oq�r�Ԝ�1���n�`	�ֻ���Q���D�g�i�͞R�H�٥b��gR� �7A��]�J�"�����Df�&��v�3x���7Ȗ��|� ��N�V�Uݶ�",�,�=u�a�T�M��Qė���A8G����ρ)/�����%��Qcp4/��:w�v����O2�!\|���
��c�MF,[v�Iػg9Qu�;|�2���x�ee��>f-�����v���4�B��[ia+�?�;��If����p�Q�Df���Q,^�R���E�@7�!�5�W�"�C��~v�k����>�S�O^������Ƌb�D��,�;���|��H���e�g�*��IS�Շ���N�K��R rWt5���T@������H��g�猟V�n�3�N��1�$>���X��a"38�<���/=ds���s�P���3CЁ�� ���`fJ3~f�x��L}����8��`�d���W,#kX~G�'��c��Hb{8��Q5��n�L��h�L��&㖈�y��Z��Ps+����J��q��0АO�e�s��\g�m-k���Ӷ~ৃ%�͚g�U�\���=�b&Cph	$�z�.I8]�/�����$/�
>e-TN�����Q�K�X� �CL�����ȋ1��e�Y%��Ф?*�)P��6H�Ì-�X�uaAZ�RM�5��E�����Ill-�cEq��t�]�'$�?`^���(*�A6��8Hiy9\嗨i*�/��TT7��M��+� s�SP:���;���$��I��a[�lw�D]��|���M����f}t��I�*au�A�R��Z�uHЅ��ekEvb(i��f�F��xx��R@�oO1	�h�>��n��"�M��'�`%���w\եT���.�G�u9S�Q>�u��/f�_"Inz�!�e S�G&q-lEe��!�|K;�VO���Gc�pQu���M]Â�*��[�>h_@6�v=��Rf�>ʯ?9���񹰐$�$dV[_�9�,��l��7�;�b�T�T��f�/K�!Cg��b/��D��b�h�#�q�n�oq��R�̝dj������FNd)H���p����XyFL4�x_#jG�̪d�	�	5�S�*�G�.P΅����p��2�Mj�i�G�0���2�f58�Q�I��ܱ`�fC3���
�f�#
3_�� ��u*t3E�sd���D�ϩg�g'�����c#,��D�P=�	���S�/�o�W1^8w��b�=[DO
���c�:�o����=�y�V�T6s�pQ|���ItHS�8���GI�CJ"�P����]���X��{�ig�Ôf���6�F��1P*i��3��\�O� �.�.)��J�|o��A���k�B����\�H�F�����`RLZ���R�`)r�j��B#���G:��0Jv��^l����Vr�����Щ��"L�1 W��^��Pd���;x�8�d\�+Ly����+�3!u��Քl�h:�:}��=:S��T���ө�r��bXc�Lګع���=�~����CҾ%C�e�'�t&��c�^R��bSd`��M+���٭��#�	����&^�NiͳP��e��Y�i�&������Ě������?aɗP:a�L��uY�L`�t1������o[(:�@MS�d7�@���A�gD��#��:L�x���F"�<�V���^��a�O}��Z��:_��7x�Yw�N�ަigpo8�0( d����#��^�L��C;�9��5���.3�Wi9}�lC���y)��#z3�����3[���$�@+'�����n-җF1��CN�Dz�ڒ��n����hd0%�wlM/e �\中����'���g�u?)7��e������(:�h�P�]`u�Mb�"2����8)o�ohKwdI�b��V�ȹ���Q�u��������?Ńrx��p �1�.d���թl�2�T��)�K�̈/�2�W�~"�Ru�6��B%2Z�^d/i�#��U���ͳ#cj�S����?�|/h?���+��w%��$'!��.]֟����ʆ�8מ�X��܅o~�N=�:,�4��~��%�F�ch��:�4r�$*�N��l� ���.�w�RW8���`�.��o�$��dFiVzR{����ᎃ[�VTTka畸�1)֙}��o��G���h8#��G��.�7)X�ۓ/���0�����AԳ����Q�%�VD�f�{��$:rM�x��TR��?{�������#��R?��p�m>}��شwx���νU�{1O�ǐ~�Hx��xX��v� �fs�z�i�?Dfq�aO9�fmzu��
�R�(�Vmv�I��;��U�p ��\,���|Vd��Yߩ���Ρ/���_2� p{}���I0�4�V/h� 8$��7u�]mL"�:a�:��GHE��١/l���f���cEɎ�U�UJbK��+�R��G�O�+2���Q숸	z�'7��d���F����,�����7���M���  �z'k]�������ϭ1u䣊���B�Ǉ!S܍��.3Ra�O�h}{�����T�6�@bŢD�X�ؔ�R�l� �Nҩul���Ƣ̅5�d��H����D񁱵M�%�ӎ�l[ʈ C�v�,*�g]���'u8ѣ��{_m���b�{�)L*�uݾ��1+�9��	i�=��ۼ����ɸ����M[VS��T�n�����OG1CM�:�Qt��(�ѥ�j�Ļ�A�̀�ӓ>u�1cEM�{:���i�PDtX>"%V��}L'��Z�q�l�+:���×�*9J7)N����ѻ,��
����k�����E3J�8Ed��f@�H�.�mG�0v��DS+�Zp����Ӟ�^���<�N�:�)��
r��6]!���/G"��q�Zp<?�_���.(z��# M����z]^8�b&��K�&#ype;�����]a�01�`˙YdN�f�xhC��;������F��d�OE�ǐ0�,;&^�P�4cK��� e 
&��ms�o��7q��l9r�!�)�f�_[M�:��SB#��Aׂ<ʃ��;cBv����@��ԇ�7�lG?��ʤ��� �U:l�\Z�&|X+z{�z��a�SF�M�A�t��8��2��a4��נtWh���;C�xc�����b�x��eWY_]�Fb�0Nߢ����㋞g�.2�х��t��>1�ƚj$���9�դ� �6x[��1eR�}y�  ���CS��V�0��۲���/R�N]��Q����NO(n@�m����̞���ɩ������&=�*^�?�,[F�	��vM��QI񯳑�����Й�n#e�
z�hq
V��f�sTo)ո|�Ig�@+�JA�I�}���U-�Ȅ���>�<J}�p� �0-��U׆��y��K����/��[�ag4T��lA�9�H
�+���nĪ�l�U�L$V���bܥ�EQ��9���8�"'�a	�� 8u���6K�l5O�ڜ�ڜq�w�e'���&e��9Ks��o�1�����G��ùd:����ɬO�Sh"R������S}�
�^*_�D����������"�D�`	! ʎD�*la,��I�q� b���Au��q*˗�82��gN�=��zW(��ф��X���0䅈�
Q2ns����y�͊��� y���z���Mq?�Q��0l_-���8��1%]���d�Y��UV��gV1ׇ�J����mJI�N��B��U#�u$ύ~5>�YKQ�M�E�/h���T]m6B|b��1��PJ�Mڻ&cZ�PE�]o~�*�1���~���N�������8�����T �	/�qQj,l!E�qK����B�˨ |J�����d]��Ìe.�p����U\
5�]�{\���N֎]�t�@49
u��ǒ�U��� [Gm(G�����KHg�(��9�g�}��R@���㎂� H�->�K��s�������  ��v/KD����1�F欰e7���T�ɟ<�2,RC Һ�扴S��GO�`1�Ӆ�v'���0��·��%��-2`"6��ԁ�c���q����[�1�u�h��x�ƺʳ�b��A?fODh[Mf��m�'�:��>�;5y�v��PX�u���}���^<�f���{�3���9㥫�ۄ5��d*L�)���A=l��#$��&\)
�	��cz�m�:Q��G{b0�3�u�s��M�-��Y�4�w\��45��R)Mԋ�M�����$��}$b���>vd�{�'��	rIY��2���4Ԙ�-Co������W��<Yj��)�"��:�
9,/ 	��)˅�h����A;���N��1p����N(��4�O.@�����G�g�s+f�[����=\�
ǲQ��"s�zv��%���z�>/��0�f{�
�<�+r,�2ښ��K�W�䦻 /�\8�X������]x�юw�%P8��Q�^����ou�|v	�4�ATS*�z��9���4%/�[�*�/�g�*'״@!R��m���"���X���v�c���F�-B��Ou)�1�%���/��)ӥ9��6���TR��B�;�\m�;� �>�t�^�����k��3��G`��t����[a����=���t>8��J��DF(<r����F����	a�!�����t)�tl*�0��Q���WZFMf�[���
�$E����6�?M���Vs�Z}�d�s��03���9(�����/	�2�A������Cs�Ȍn?�+��yw��{�������`M 
oe,��=�+?�y\Љ56E��ϖLZV�~�X�����r��C~�eTreD$[��߁��a_`�!Z�=�9�jtY�ߎ1m��m)�ti4)���c�`�H���E����6|���J������P��5�C�m�+��bq=C��y�<�$e�ibѐ��t��V�I�c2�VҀ=G&�����9�RX��: 	����������!i����Z1�C3����e7��x�e	��Ѣ��^O׏��))=�'���
u�N������#��ߩ�,���?6� ��k����u�8n��*�R�l�2��S���yU�٢�-�^W��az�z$^&���1V��&�<��"�r}p��Ճ��w��2���c�����cm>V*�r՚�Л���˙Gh��ƀ"W��5��d]:3+9���dF��V\���>nW11��=��G��1��u��omr���1�,�V�����5!�[1���=E2�IPʺG�<��q��NxK޲���a@ȁܦ��0 C�wAUH����$Ȏ"`6Vfqⶸ1-!�G��yQ,�W8"�hB$k�������}��;�
(�L���WB�J�FX�ѵ���l@Zϓ�_��)vX�a_n[���Y�@x��(���F�!K�@|���m�m�P/�n8'�� E�B�D��|j���.����2rhˎi_�xM���E,3&�2�����u*/���������ʚI� )�N���(oy��)��HeI����I��ie$S��>��Iڲ|)�Q� ]]�1?�ُԳ��أ^���9	\�++���J�w��,7a�
ƹE)Z��K@�=�D��r���k/S"����Õ�JQ��p�K�q&d�I�h�)�Z%j,�9��ZN�#d��(r&���{k�M�9�ʀo�����A>��3�I;��!9s��9ֵ��Ə�3�J���B��k�!�.��|J��#�S%ta�z�P��呸��_��tC��M�<P�/��F�mVtL��0���1�s�98dz�H�Fzn�����)V��(����{8n�K�$"�cyvD�n�Z�h��=�բibɖ�\���Xٛ�`��m	x� ���T��d�����6<H;�����6��
fbx�^�zB���zwW|js���՘a�ӄq%� u��|�W-�X�YU2���Dm����s���jrY<���;�|{��_T��%��|U9_���� �J� o��/�����O��zTƁL|���~�����_��1�$��Q\Uz9�"�{-��38֑�TI���T���.�ב�������R�9�M^d�Kƺ�D��*�!O���.c����vY>j��'=�>i!^\cg8�	/�@i2ݼ}C��R��*���	0A������l�qA&��ܻp�J�"z7>pk89����zq��J|���w 8&UB�iԫ���mʔ(��z8h;�VB]������%��y��*İ\@���F��5���бw�U=XPV� ��ӔaFu�Pu�[���xÀ�B%��s
�-�V��Br��icB�}�j1��%�/?	lf<���n��4o�}�����b�tP�q{&}F[a���Bه�*�<�&ɟ��pjT[�%�KK6jQ*��W�KW��>]���l��c���������G�}����vv��6�ru Ou��fG�kExS���!.�o�֧t������\���"c&��� ÝY?�M /^�L����a9��۶��Y��j^�����~=��R�o�ZOY�Ӗ3(���;�x2���-�!bD`N��/D-��n:H�9O���7o$!K������]e�L�����9��%�*%q��A~�R����*��N��T�K;���*lC����K�@7�/K��R���R�:8n_�e�U���A�-�F/��*�!~��R�һ�����XI|�o�� �V{�9ssYQ[ǟ�d��<\Y3࿉ْ��[���RZ����`�T'���X7mo�=��5[֓v�
�;ߟ�6�e��<�mw���켓l���%Y~N\��^���/}��忢s+3�S� �Ѝ���1�i>/�q��V���\���П�R/��+c	�7N�SB�0,^������������v�3�$���t�q�� ɶ�ϸ��w
�Xŧ�&'6(�����Ӽ���#-0�d���o�0�,��!��7�l�_��oI@�n���yL��4�(�#�L@O����x���t�+�8���6�'�p�$c�ЈQ��;C�O�p���>�B����V}�c��[�Y���$�B�J�4,8�mo���;��B?�|_$�}�C�*�X��a�2&��ubɼ6��9,Ta5H�5=��3Q$dV_��y��΅Ȱ�[�N��.��DF�Р�6� g	!FW�Xŉ��o���ߘ`�wY�f�ɑ��_��'X$J���O�6�������8������P?߇b�?��1`K��̘  W�0�|�>n�*x�5�sZl|5��@Ç�D�,����P]?���{�v�6Z��N��������<��#����U�(�i��L�㶫�9���`�#��4Y�&H��Q5Â�_���s[��V�+����{�A���'P7��򶟲�1뇏Cd��M"3�4�i���FD�:E�K�g�@|3��\�c����O�]���\B��dP�C�/�q+�]�"�����y>���6�{f�q���o�)�l�=;yJɀ�A�z�'�뀉�/7}$
���m?��9��2Q+��l������(����&����I ~_��y-;G{j���Te��'�˙XN<(&����JdҊ�Y9�������y7t���mj��bM���rE1[n.�1/xm�mA�0�h�pc�ѾOz-�C�D���`��c���2���`B+� -�Pp��,ǡ�]#[�N
l��S~9�!qZ\�M��� ��:^e/�\E�i>�'>M_C��ۆ� I��	<���3H��t�������iovܐ� [����0m�2����v�����,[�w� �K��*��0�?Tv�������d��z��S�3wШ�����/�6��_�)����!������Jw7��Aa[�p��"���}U���jZ��m$��_���1
J��,u��#wy~��~B�t�`�d�?hh����ز8n)쌖����3?�C�d	#������z_1��h��MUW,
���-����rW�b>C�:�é���~X1��N]69�I�[�!f�Z+��������x�`v.���-6�4��U�'�����fA](e��6�T��v��R��)�~ȭ�04�J�NlNG��!����`���b�Ӟ䬈n�O�3&�+�{u����C�R^|%�j'�yE��m�&�]�.2��j&�A{��ə����V�e�7��8�.\e��{�&`�6f�{,C�Ca��fݼ����R>���m� ���mF��m��TO��#�5��>��[��(y�4��[r�1�t.���4�'F��&huU�������;���^�űH� о!�`K�yOt�҉�1�ڳ�u�j�����_EZ�Ŋ����H�%p�2f'� ��0�d���LS7��=/q�e��h�Õ<�[!!oe�@��d;Ѵ��&=8�tJ���f�\�q�����k������VUp��э0R�o���/�;팖��v$LW�|dH����!�Ӟ�x	goԋBe�y���B�R{��m����%�S�n߰D���Eٴ*b�֙G�
�EP�P����\N�I�"b��7�EM ��~ܢ �ʏ�W��u(�)Q�[%v��;f��u��y.2���I�G���Ry?A3�U)9��m٫F����kH�R�r�'��
��o͔��}]��ն�4f��u����ʰ�����l8<���(r��\�\��%����\�U��B�&ٽ㼈�y _W˅Vq���zr���ȼS�3�iū�#��천mH�B����� ��H��f�F�2����'�'4D�;[��s9 *���	�1�&�������1HPd��*�&�zN8�c��c���b
��:�࿸��z��kb{��=���W՟��2�W�����쬡�$�]���K�O��!S���(%�|���^U]��`��|_�nT���$�2m��y�
M�|��'�BNj��_�Օ�|����g��[W�ї�����#����sR�VT&a�fp�>W�is��wM���g�i���ra¶d� kD��ܽ���Ƀ��?*�2O�	j!:H���Či�Bݟ�ᗬ�~"�C��, 2S�_ ��g\R�S�}m*7�󖻢MY��Ԣ���y����;�g�51H��t�Y�؊Əޭ���d�C�p�[�����D�3����KB���/�+ՋX�o챁����C��I�|�f�-XT+OIw��*���p9��g�� b>��b����{F1RU��N� @K,���$_,V{e�,�^'�3�]�P2��bK;� i���?9��t+�F�'#����/eF��`X���A�N�~o������5�.�$I�E��%�~���ɐ[t�h����4��;����|gҎ�Q�q�e��d(���^�p1I�Z���V��*��4�[���򑮡)��A�����K��Q��RTU�(B�g��7N[��X�E����	�W�k��J"�c�𺓲`��N�`��@���t:����UB��^<�A�ȑ�PD�VW_q�H�g!,c�^����b����i�j��\���c��SB��MY�r7)���U�m\��?�RS�#�wW*�e�Fg�<|vCwؐ�;_��\rOc�|���D,8�B��v
���g@v��F��Ĝ��{l�ء��_��R���o�'�:� �\�#t����z���YY�
�1 �2���`������$�bv�g0`Wj�����y�.�ߐ��@E��%g�#\$��s
�?9��UPpƔL��`dK���j�����o�p.pE��[�jU����MY9�G��,�4n/(z}_�h�H�%��:|gm&����1<{xn`����Χ>�v_6v$��i���%m$�{���laP/D#����g��|��H}a���_?���&���bMeTK�w����Ү�tS�bKδ�ʗ�Z�D�u-ȑ�P�D� ����L$�:�/�l��Z
���D�*$7dQ����6.�m����݇�ќ��$	�,k8b�����:�#J��s�.V���SǪװ-I@5�5s���j�Y-��
sԸ���h��F(����lpҀ�ښ����в7������d�D�{ڸ�$�C�Հ��T�i���`]gRQ��ĔѸ�M��٥�۠O����J�w5��YR4���	Rm��*�I��p��D-N�sSj(��E4�Md#��^���d֠s�:-���S?���������9�t�A:�_��&������Km<��ާy��tT�*ݔ��L� ��V��"GF��F��	��2����.Oo^��)ջc��{���9w.w/�M^t�?�Q���b���?e2|׏O�[�>:���'���>+�n'�ࠂ>�l~�����%���yfq����j�2?�{�:C�q�b(��<�s��`ǀ��Ȓ�Q��~o���gm�籉)�%N�܁�YT��Cɥr�]�,<A���M_)�ӓ�۰�b����u���8��~�W�0�N$�߮O3d𵏠���tYց�i���r~�k��?6�W��%sV|Ӈ�8dc��G�*������?Z���P�d��0J�}$���Vyq��vIa�r1��͌�KJ0&�K7y�����Dua�؁���cx����=���G�@;�M/j�	���������0�T(k׼��'��`/W������{���3�A����zK>����f}�2ms��ש.�`����deb9  `w���`��ex���7��1�R
�֢�sƄ������f�Xj� ��.�|�@���]�GLp�s�=+�:�섟��o�Dy�^�+A�d4K����r������(Ld�6.䩃�G<��D�ث�;E���evH�3 �,W�ʌd�X+?8U6�g W�Ż#pʓι8��#��4����vO���Mm�K�n"� �o��[���7�:対B�(m��b�\GJ	hs���&w.�0�:��|I�_����,���J�
D�F���ڔ`�Ȝ������Y�v	��7����_�o�]-�2���y�����N.SB&&����ꓟo��g�K�<"��� s�YGL�����1*�{�����)�#��.�D֙y1i�kB��R�c�������A�Q$^eNW_�t��g��[,���t�_�%��^..���Hj#���ٖ���{���a-�ʦ�����`v�c�e�_˽Cx��n�@t�}شQs��ڪ��?��!�N�w_����6�<�������ЩY���i]�%�T=���/_��*(�sq��l;`��� m�cdtv���&�p}	r�'���"�O����)}��_NM:��_����Ÿ��a���M��Χ\E����׺rn�2%��S ����(tC$JO�>R��dGG���YE�c��U��tZ{�I?�D�0�t�kN�l�$&F@n�5���t�Ǌ4�d��4���>���ǃ0&�;�����g�=�,C�����B��i?л;O�V�m|�i����j�A��*��ZX�7��-�*��[�b1��~kZ���B(J1��K0^g��F�C�son�,�3� 6��u��ͧu�._qWa�����]�N�XGR'�B`�t�q[,.+'�o�O����q�����Mq1��F��������vj��K�Gɐ O�UEU;Y׉��Y�����z�	���2��Cl��؅���p��aё��|��]3�4�	�z963��G��QD�nuAU�W�W�j|�C�
�Uz�6�T�u=� ���Bd�8}:NV��Ɓ���u�#T$��}���"%�I�=إ>߳xk,��kD�(-�X�*����B_����M�f4ո��P.�B���m�ۇ;��	Lp*��zr>�E�>�GŲ?Ve͜-;�c4������Cݳ�����̓Է7+?��2��6D�c����I�\�G�؞Yr��tϮ�i闰^��U(�{���.�@��U�} ��w7r�*N�n��8Y�N��q�rٽ�M���R�q��c1�h��]���Ta������ʻ32m��䛝t%���,�t>҉6��m�9&F��`���
l�iI��%@_��]W{��a���a�q�H��Z��VEΆP��U�?�V���t7Goj@�$9�K�+	��[��d?#~�{����OpS��������h�g� ��;V��_6���8b�X�탨yG�����?H��L��!K��*�C ��T��U���<J� h���K�&��{�+��΍�R�\s���+����	G9��C6o,)��%�����\���<Iv�e�z�\�G�J�'�#=�{��ן��H�@I����1!F&�,��洸7	z��, _Ȇ��Z+:G�ѽ�,$�V<2E�ٳ�-��"�%G �P�s�W���l0��ӝ��#�(���7��$|����I��pK�⤣x��Q�\�\��I8��/��^E�q����o('����d�a�[�����xK���1+�{x������4јu��)�U�x��O1=:.� �"�=�g�aA��KlĄ��B�|(Aqn�N�Ǩ��yh��8�%�������K7����K��}�af�Q�Ștk�~^r�
'��Į�&�t�U�m%e��ʅ/.[f�j��>U0��͸5��OH��&쒑Q�����`�,��.0��׎:茔k�v§r�[���F*���;f�xx$��6h�U���︒�,�@2���y:3.��i6�p�W���,5_d[xډW1��1g�bcq$G��O9�8�^�t���N��� M1W_m;�l�Ox/w�D}C �G����_!��1j�e����z���#-k�����(�kt~KԶ�НB-�.̛�g�}|�B�Me���01��b�ͦ; �5)��='�����3&�%ػ�7����JT}�˺\���>��2Dcl��gi��>/̾)Y�Vt�¾��w�s2��ֆ+�q�qz�[U�����m�8��gmaO�n����+Tkk)���n>t�'�[�8�����7��9�  �6#�9�d��
z�\�Eһe�����oKٸgv~�,n _�m�w4���t�}�;5�佫;�"�8���(��޻�%�9e`F�_J8��u������?`1h��3M�B�Չ��6���Y�|k�G/�`�J((.����I멖U��z����A���do:/��x�:���^�������w�ޑwB������\������/��X�����H�ʏjZ��9�.�t.v��d�~iЦ�k�M���X�j�oy� �Ϻ�/��x�:d����擞�^h�gĢ#XE0o<�q�Z��5K�{ԓj�>t��
��L�k��#pq�W=�.f �~��$�0El ���ì�g�L�?|�.Z�x����e+WǠ���$L�G�7EZ�V��s�A��8�X�d,��L\:y��?���9(t������t��u�d�R��E4؄U6�����-���ȴ�O��qf��WY�V�Uph�n�e{1��%��< �Ү�]u'��SGa����[vȜ~X=-����>)q��B4�۫ �T��!���5O�r��.P[/RSHW���B&�5���yL��