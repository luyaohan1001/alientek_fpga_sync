��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��zW�&��dO��!Q�����o�r��ڏ���U�Ta�T�j��\�I��_��Z
{u�7�S&b��[QLmP�٩��	���'��>4�q�Z<*Ýg0����8���jܠK)o��i���E��J�_�9�L��~��p�9zW�r�ɀ��0cUR��:d۫h��h���tYzT�v?%#$�pA�%:F
�? ~�\�S���i�|Lp����PMd�'�a���8�-G��1"j�(��|�~;�BX
�x��!�1k��B�I�����4�����P�ױ��Z�GM̡(��$�-�4��
7<n��%D��0E��0�Ȟ��9)������G�r$�!tL`.yT����AC4�I��k��G
���A�i��M��z���Von�f�C��.�X�
�|�^a#c���HhY9)x"ٗϜ�����p$�]��>�[�����ê�tg�ۇ��v7��O��|�H�L�����)�{�I4��N��m�P���r��o��i��Mx:�F!+8JVfX��������%4Hb�+�s��漻��rf�*�JŜp�(�5*J`���ɻ;縊��$,5R"�<ow��%5B��cоK��%��Єt��/&��+�A��8�l��*�7)��}��&(}�V�R��;�E�k��k�E������wA�K0��#�yɱ���`��롙aKz}��B+�%��	S����E���T2�����̀h4���>ʛ+SG��-�E������}�݌w%��z�Q�qGT�{��i�����nճ��T��3��-� 	��s~n3����;j��V/I��q'C>���D6\5�u�y$gxo)o�C�qT��o�%J��V���ރ>N�8e���ޢ���\���(d��|M��pR���~�
܁\ɶOS�]�8�	�' ���X��[�
a���S�I]t��2ˡ��,�O����yJ~f-��=ק}���-"�&�UB�ܳP:����ji�룣]����F5�wS��� �uױT�^F<����{�Pb-���j4�y����8*�,x-#��&�]�*��1����O�l2���F��]昹3����^)$#A����mF�V�k`Uw�x�(���Z�Gg�5^&���xg ���z���'G/�ɮ�7����}��[R���_�0
ƞS:lv�o|Em^��̖l�"����^�2G�ͫ9�s���"Ѿd�$}1�0��?��
k�ǈ}7Y����2�_�����Oo��*L�2Á��ʶ�^�O�LʷY�u��c����n��2�|�z���IGg�ZP���Ra P���7���r�<(~9���< ��S�I1V�B-�l���5�P��$�[f��ph4�(�0\}�6�`�`v�8U�qq�w��h�NƓ�5���,��IɪHV?$���Z���&G��D��35���*����G�N1����#���QS|3������C(��ժA���r�F��;�La
˗����6�����_�ː�3��)��[���7�ë�����`�z !��E�h���I(!Pi�0& ݖF����m>'o��ɒ#�ub��o��%`��.�C�i�9
�i��!�pu�]���)RO+8�f��m����Q[#n+ߥ��������9"��9�E�i����t�;���ɛG|*1����MeG��n�z��lrJ�?m�0�'�Hwg\�Ɔ���_���ϻ�g���=G(��9�N�������j��L�X�%ᰧ*I'�p��o�vB|�t�Um��܏�X's�LC\�%��'�AF �ʲV�����d��#AAx`s�������!O�*�} ��!V�	h�؂��6�{F�[Ay;"k"���/���[9δ>���ڪ�kmt�{,2cEx�_ f����s�k��{���g�{���ڀ�PN�_�kG��_vΏ�S�	o�R�j�3�*�ˤ�'_^���ԡb^B�J7ҡ��K�a!���{��I�h��Ȭ?L��"=�� �Nh����c!t!�-�z��U�<h�	�0��f��~G��!�L��`,������j�o4��3�y�V}ͷ�� ��ǰmɎ��zĲ��t�z]��sZ��1� ������đ�0"'�HN�rP;6�$��_�vb�D�I�3�����'���F��Is߀�X���W�U�W�:JŐxT{\,�u�������:��1W��P�\�#{�i��_���-��M}],𺒰���d��, ����KԺ�WL�ǂ咏�<h�-��as)�P�M�.�k�K�����A���Y4��T۸e�����=��`�n¨kK/Z��_6�09"���4���̰�п��A��f�m��U���-vZ��[�O]�L����~�Zy�
���\]��[w�;q�Z�S\�P�+B���N<��sUȺ[�Q0>Mv����#��Ĥ;����g�P���ܦ�]2ɟ��H��ףÃ�Ⱦj�l~�Zt�p�)E*�{��"٣����A���dC�Oo����z9@�F�������U�9�SI� ��Je9 :���j{��^_N��ӎ������YC�+�B��a�m*u\6%�F��:�0:�$7z���c��ip������$�ߡ�P����2mW^���߁գg��1�ac�蘫�NAO�+[
`�b$�a�1O�d:�X������]��M��%�:�*�?���t'���8��_8I@��]v��_��Xk#-�q��`�x� $lT�(d~k<JIa��R@�?� ni��������9�{�~������Wg�8�,�h.��`2	Ae��/�e���FDAeW&�c�MW5���ϙ�<H��$0X��M��^�}.O���s��X��Ϋ�%I�b{�\ʽ���b�C�Q�8q_�_
���&w�g2��րxT����n�,Dra%�+�2��0�����q@����_}�vA.�8��ã[�ڇ�"\uCO�1ⶅK���ng3�2즣�ě�]�k� ��ʲ؝G�ջ��VR�ᒡF�j������l;w�Y�Mo��Ta̻�
=s���Z3i$i�?ǝ��d���v�x��T�k����N�4�<��˶F��5r嬭���jek�6eH�KC���4t���H�<��`dѦH�bD5F�]�eoڐ�O�1��� �����"�n^q����{8|,���5�!�^���y!�ңN��ao��H��j�92]28D}j�/*I�uy���S�,k������G�k��cK>d;�z1�lj�g��@d���`�/HQ���<�'Q�b�}�� 4��b�r�$�W!�I��œ��f y8J����謪�i��thA�WF0=Rٲ��	�I�e�A��lq	�k��~��O�>��Y�G����ޔr����y@[��,}�W&�*k0� w}a<5fʛMu����>n���/H�������*
8[�� v�U�~��:,���pV ���d���-����DZ��Y��|az �W��%��	��`������.V�6���x����$hg.`�A�[�`=���U^`��y�z��^�w��k���ܗ�s޳M�>����C	�6�o��^�nersA (�Sԯ��ʅ����ò�Xт��ۓ��"V�c��X����j�Φw�f5���8C��zL���OՉVй�/�|�O%$A��r�O�gI�ܔ����&F�	>��xz��Ki�<�x��c
,���naŰ}�/����E,�i������S��W�ejw!��i�g���>�u�w`��	ՇY���s�}ڳ�;ִ��"�VM�p߈��BZ>������`���sjV|Q�vL�-��!t؟TCnKFvҚ寊� Iѫ�9���-FSuU������T��kv/��A"�RI�(�C�T��n�����YB$���/W�v&2���5% �%5�{l8�Ҕ�'�d�H0]RɴlZ�~*��V/��Y��Z*&�'�H�*�=j��vv�M�Ǜp;_%u z�l������n��P%�XzBC]�̊<D�H��t���ޤl��UuV�]��e�m�C�!_F�������r��5�3�
��3CAh{��v�
�2�:׹�Pd�8G%|�"d�ر洍���g�ռQ��L5�!���(l"^�.�"}z����4,��v�{	�0�6�r�y���f�+:��C��ڜ'iװ��0S���Eۨ+V�Ơ���R�J�,~�y>�pW���Fxu7pw �k�����L�m�W�*��s��l_�׻7�[����h�Gv:DY���=�s۵>ph��G�Jšf���!iB�5g��Ud�W����nb���
���/ ���Áb�Ѿ�X�DlJ�?,��x�j��&`@��t�p�I���ʇ�"�`�6�s];*�D�ǂojW����\p�I")U�=B�R�,�6��m�X��@U�_������ g�0"&W-^1ߨ�jC	8/��\kԲd\^_o6�)���ΰq��M1���d?�k��������ߔ���C�;t�%#��Hb�\[�_\3�� ؝ϗ��p����'�F�5W�1%)j#�@%Ku �q;/fh���R
���D[T�?L�:���Tpr0/�J~��'�&��5F3 S��>@�5�(���Qc�}�u΅%�_"�mπ��uw{��b1�j����w���[�����>�
zO��m��Y~���,�����5gt*��S�����H��b�<}z��*�s����VY����j<�* Qd��ɟ�k��tZ��_�����up�Q��~���/ �eY��X44hՉ��K�������1�Q��#.k�שo�V�c�$y��e�ҽ�=�ݹg��j��>/3���ϽpǞv�"��,�@��_~F��74��5��?�w b�.}��s"�oq׀=F�?�(ކ\���2�:hi�3��+ز������A���NE�T���$�}�Y��C�	�����-`�Д�X#Ч8�=ш��`2ma���z �-�x�Ej��"(���*ԤGpM��?���V �Vٜfw����[C3+r�q���/�f�<��T8�C2��ޟ��~&�/����8ަ���s�1�#���ݣ�Q~C���{�@�0�L�����I�"�>�_7�1����f��~#^5N����@R�C	�5����'�i7C!��@`�ރ�ڦ !�5�dF��Q�\�E�Ct�N�e`��}�C�Fz!p���˅':�O��B�EUח�W�9=$�\c�(�FeJ�	�e^��Ws��9\Rx�Q|�����g���t�*(Z��,�~�u��
�F�����)��,_<���d�q[��jE��-�D�~����y�,:��Z*���l$	[�L�e��B���g]=0�����t�����q�w��˨o9�5MX �0�������N<6��p��� �l�G��zU2��)�!�bIĺ�	| e��Њ&	k��
Z�������]q{��3�ɕ_�����6�B�h�L��8�8S����2-Ϙ�:�%���a�o��:;��6�b:Y,X���p�A�8�h��J�94��M 9ހӮ?��ڵM9gbm��)#��H�	��2�ssT6D=�n4�%'�GQL�;�xW!��O�I�#UL7{��b��Y9(�V2:�=��6')�U��iOl��Y�v`�:KkF�Қ��IC
�63�g��3�4,ڀԢ�N�Z�]�PG\ʣ�꧋�킓.UCzm���m����c(��Ϡ83�%(7�����N�CK�4�I�1��B��l��Tz�"q�o���B�tSM^sw���hw{�j�J�+ ���p�\QEu�	���9o�u�Z�Cp�4��A����o`�O?�)=���~��l-���J�9	�R\?��~� Lw!��
�H�6������:Z5�_� <l"�|���IP
���0�v'D���)FT�p����(^����ؚ@��}�PZ���'�����M��ڇ�q�ƀ�ɴ�������l�����݄;9L��β��ǎ�WhC�f&���ù�Q
⟠��o�S�߱�8���Wн35�B./	rM�H���cˉ
=%я�J�Nj�ج�+��W��q������c��5<�a���E ��\�nfL���{|�T~��������]c�gF'����%��v��]�B��ʥ/��� ZM#.�� U(@@��n玱#�0P1�"�"۶p�����2�!�Y��}�gM(�靳�����	��<
v/���Ƴ�M� �ҷ�6�y�Ij̸8�֝�&焛�����L}�?N�Ù��b���л��s���Ͼ�H;��譐���y�Jg0��c*��˟���!���z�Y�����U��MYĮ��l���<G�E�ne+Z��E�B�~9M��T ڝ��Y�$o�^����<F�!�������<Ⴑ<iAR,R��H�I����N$������)��dk��`�&[~��{A�i����0Sף�81��6�-�eT���+(��u� �?ڋ�,����3��6��_��.5��%�k���x�&mM�
�1��w!�?��F�:��zz��|����������7�y}?8*!�!���L�V5p��ȱz�ɿ�t��e&C�l�׮��[�
yYWa[��n
��|.��i�ӱ!�"�Q���e��t,��*O�0��j�d��@�B��o�G���1���dJ���u_��E ᆵ���9�1+*�6�?]&Ɛ����"4��_`�oV�ƞ��O��QJf�z���#dꢒ���%W[�Yu����Bjd���߈�F���x���6O�~N����;�����󱊴�"<G��5f�����=���9���BZ�8����L����_y-�޶E�Ȇ9cs��}Y0in�I�ӪϚ�c�oPw� 9m7�%8�$��&��g*J��ho.�qWx̘�\@�͢��xa���\� ��h8�'m��iQF�OF��	�믓Y 8S����Oz%2�W8xw�4j�;�F-8x�	�����K��.��{��?v�D)-%|���*���F^=���͒�&*�\��xz�<o1��|M�s^[��=��އ���WrQ��
�,������K���=u��$�AǾd��cY�,Uq��V��=���6>������a��p�(8v���f�ׇW51l p�W��q�a�v������`����E��p����3P���-VL(c%��p����WT>��g���
�g@��@[��0I���WaC����Uu�w,��u�R�����X,A>�N�P�9i�0�c�H�����t�g,M��jX���b���q)b\�)K�1�����DQ��a����!+8p���|��*�u���F4�:�_z��kɃ�r���kA<hr���aPve���$y��hF�pJӡ㍔�l�[#�HV���8��'W�M���L�	*JC�#1]��&��[g52}��x	�	�YR/8D�aS��ic������
���ܰob.2u�@��J^c�O�L�SHq�Q\����r\���q�O/n�+B��Ć�{0Vc>c��d�
븐���A��p35�Mp@\"=.S�Qqfr{o�+KQ6V�g;�ܯ���ٲ�]� 	�p2gF�gI����M�"�z�(:��(��05�����6@��� ���	��!P��'27�����9h�����O ;]B��Dh�|RC���a�A� Yj���1P���,ߡ�Do��ף�z�1G�e��i�v\VM褸K+Ī�;� >i�{�qfH�Nl�Q�8?��rʬ�Ɛ)�״b�ǜ���j�����u K��L��,X���+Be�����	�	���
���s���g�e�l�(�`�`6t��ݔ��)t�D�yMSY�VNߟЌa�[*��#��[�J?���WڕW��1��j T֢@^�-
��",��h=u`�t3N��^�|��	����1%�����`	� {�G�,���F�s�z�,�JI��NNo� �0p`XXi���c�e�����R6���N̴��.!V=�$zA<OZw�Z�̜Bϋ�jfo�\4�����%�箜d��,���N#/��$V�ɑ�3Ydۇ�M��(���O,(k��qUTb_q��X�p�L�:�$Ub2�ϓ��RD��·)�L��ϙqT�a��)��E�q)����HH_#�e��֖��F�>��,zo(Ȉw�*����L��M�g�]fa�oJ~y�h�SH����e(W�(�V��]�����9�7a�� ����X�Ŷ�,f�R�f1��H��*�@ݞS�T�	�#(.S���[��Q�2�0G<䦬�Gѱ`"LӒ��6T�����%�W�0R��le����(�$���PT	Z|M�`"\��6#Q|�@L����)R[�po4jI��Q�=n9L>#��C�B"&(���f��r>WP�֠��'+�FA����3�Ժ�&Cakb-�]��Td�k�f� &�Mxc��H���\Y�;�t�U��Fؖ�6��ĒRI�}["��e�W0ЀP֒jŇ��c��˝H�K�+���%,�]���D
�$=GRMK�r�N<E���9���>62��rF���^؇7q�4�Y	�<cӸ��s�;s�Ynu͒5�بWp�2�R�b�O|c(8aղi�CK��,�4�C_r6�솗� ����A��aL)\[�������fj�c~�Z_.��^��e�+v��9����-�l:VC��>D�yil!�tN$HB�� �w��pυ(55�t%2���ϵ�#���ó^ F}9=a1�؅{���>�_��T��}%Q���
h�0��������J�|���5�#su�VZ�m׽���@[ۯD6�>C�?$��߹�����
��ϰ�&3���yH}F^J�q�.e/��@dS}�;6�Nƣ	�1�j������H��o�
iԑv�Ur4;��5��H����jsg���i���<f���tg���ܹ�b�Pnĺ	�{�?*U�lԄ}����`�dJ���El�#�P/���8�J(�_ ��]��-ዡ@jf��Pz���_ ���8���|&RP0Y�P*g���u��S�p�_�䚯9Yݢ Ć�Z*]K�(F�=�2�w��0ъW(d����b���9��@z��AXԺ��D;�����,���P�=�);�>��+�"^�?�Rl>���AO0|���F3��A����vB[*!��~l�OG	��}/5)6����:�w�:��L��3fP�<�S�Q��Z�@�7\�a�6�p�o-��"��-D��RS���jDB �$��$bEly���p���r�Z ��  y�29aJ�X��R�Jƺ�,?q�s�I&V��U���3�.{Ȫ0�F�o]�ke.%,�Y�/w�C����t��3",q2���"�@%$ ����5riB�4��X���P�el�y��#8�k]�V���U�6��h���藃hg�T��:�
�g�n(K��cq�fJ��Gƈ&�J%3&ǓQd��=UP��_k���
�N8S��>/��EBUV�Pc�r��0������^��E������%}�lY�q����>9��zY���K9�(Q ���I��\�2X��!?9��X�1���xaY&V@�����P2E}Y���kX����@�#!K�/��LW����n��yޅ�3Q����,%u8k��� ��[����0K�Y��]��^r���TTƟ𨃮r��>$�UZ,��2N�I��T�9����ʻ�����&CzQ�[���[�������@Vc�Z�I���eHD�İ��͞�O:��[r���$�[��}��h���Cqׇ��_��麀�)����R#�����.���� �j���_q�d�i ��w�wuB[�D��W�@�C������ �X�0;�n�79h��C?ڢ�8]����f�sO��,��#V(-�MKt���&Έ��<�ɼxaϘ�:(~}Ln��Auظ8�|$�:� �o=�P���l��~���-��/��	/ͯ�������~�+�-���\$�K�L�q�:a��u�2��&�&%EC��Cr9���i<Ky�M[4��lu���D:MJ�!����ݶ�q���OA%٪��o�c�<9�L@U�[�I>�~��O�����?�=s
�:�d��!�y��;	Q�ߵΟJ�.��W�9��}� D"[��n�7+��D,�����[J����w�\"�{��O1"��H��hD��d��f-�r���1£r�[Q�ӰAi���oa.�N?w�c���!��#�Š1�G�JH��=�D�Χ�h�����N�:t��2�G>�]	J�Nm�(B�~�_=�̰�Њ��݌j~��?6�٩��M��D��>AGN�~˝c�p�t�qp�ո/��w|�������ؓL���>�ՙ�I��f��o��R73�|���D�n���ݾ�]�y��`����%��>�8��UF�p=o-���*T�ddo���,�k�XR&X� �U����E�ڪ�;*l�fZ�%&��� �k�ҩ�O54㦡^�D��ctHG������6�t䐯-�aC����g�e蚑W�c�7�+Ҙ}�L5-�k����9AIN�R�\;y�^r!���(�nJ�1D��:HA�l�g�8��-9>��[5�����%��s���]⸈�"�MW�n�չL�[��z�o��X$z�`kx�p�%.SẊ��v���E�vn��>,ֆ{����E�J���{�EAW���z�����Uv�ۊ*q�i�Y��-���:V�Z�@m4C���Jo7����JY9�������M5=.MC/4��K3u� ��|��5��j&�'�MQx�}Q�݊�x���9Z�jM�a?���(@OF�_��^Z/z�bq�f�T�1�ˁ�h�7_v�§�}��=����O�/Uʢ$�G��!�>n0=���J�N{ei�0k�*��R�?�����9vʖ%a2��44���׊Ӕ(8���FN��[�u��Vլ����>���~����I�'�#u��z��Ձ�D<D�f�&:t3����7i�>����U�r�\�!����?��|3�(44�C���[�7"���!Ad��W+0�㷇�꺮���_��hH����Aȶ���~�L*��F� �ݩ���x܈��ݺ�g��N 4�z�~"�>}��K+������D��C�qD�� B"�c��/���c��A����B[�[�����kn�f����Kہ�͂�qW�B����S��9lFgb&v�F�q��n��u�8����Jg���X�qAq3S;�}q/��L�-�%�����Cτ	�Y�>e���㲭q�7�[��87_�@��[��r��n�1J�]��;��0$LC�]X�]�����1K��`�CN�wy������)� aC��{�Ĕ� ,�Q�/q�:��#N6M2U�I�al��q�2�b������Ua'��Yݲ���]"s3�D�=�%�w�h�N ��(�:�e�ع'����>A�`�]���/������n)� s�zWL�D���i\_� O�+�ľ?�l3ϞW�n��>#����?�ah�զl>�����~ߠv��g��l m�-���p�_e4�=��dd�������7I`��I���X:����~ɭ�}����آ�'P�6���4򹮋��������E�ߪJt�bLn0��r(�����+o=��n��j��z6���⻗�WV`���1L���o:�osd�)�E�n(9/�5霣�hϴ8�N��e~g.뿢y��ќ)s�^��<�`>>+�`8��2Z�������,U��g����4�T^�׭�c$�|㗫.���H��@��)=������*T�w� �"[rw!���f_ļ��pb���t�G�?�^�$�Yw���ԭ��y�(�X<�*|
��hd�w1\ |�M'�����[�O�f�(b���OE1����/?�P�����������nI�o}�\�1��M�A��,=hZ���(\=jKoeѻ��J�^3McDL!}\������8sx�}�sK�1��Y���U���s�X<Q�{w�q��U٣OyS\���	�ac`�(�	Z��[�Z�n��AS1�xD�G��Z��a�G��I`v8����G�������3F�XwGD<�O�Y��3�#FI�մ%#վr����,��K�=AG%�!�׉�p��M������������elW u!��(L|�h�]��/�i3Fd^� {4����[��Ϧ�EA�A�z5�,�5g߮c����%#� r�i��]\�����K?�Δ?\#��X����1nwP�
�T��g�[�12HM��80�h݈��{�t���6��@��1�������ը���Mi��(b����T�2�^�̱�?�E%eo<����!����l&@��psw�6|�q�^�q�1h�]�A�$B�6WD@
2�s)O��ׯ{�f3��ì���0.�+���g�l5|p����3c�l���V��DxV����e�X�d^���ԥ�_��R~�磌�>3k�T�J���kr�?�C �S��b��2�o�4z����͔��/��Z�!P��S�O�2��_��{w�%��˴��C�?QXh�en��3�����+؁�-e�*"ʎ�:�"BCl�����o���p-y��̎H�i"�.��|��'YǉyҶ�q���#����@m��?R�]�`���6,���������D&��E!�(��X�D���#YV�k�U�&8:��2�6��&m$nk���ɇW�z�E�.�*��̣���_�5�L�� Lx�㼪��B����p��$��0g�M 晽��]��'0Xȏ6����
��ǅ�Rt�W��h�<�3�.�NzwdP�s�ï��x}�����Xl ��3���\�齒	��@ѳL��Y�v�C`�aꍤ� �&![��Qh���0^i˃��L�1�T����|b!͐��-��	�i^��<K��ѤW�}��#!F®�Ȣl|$�E��ﰞ7P���4j�zݍ�J��&Q�������.g���Y.�֘�T�Fl��ĊO3��d�jt�{d"+�s�j����� �U���0�<�2�<��5�$q^��y�KK��e�*��@�ĳ���A�LQ�-T������x�J�wB_��������~�&]�C__����yɛv��p��UY=��2P�5�f|D��;n��&/Z��1o�&�V�֦�*�3zٕ�k���������w]ڱڙ���*/Do5#%j��-���sɽ�;�8��h��&�鯵�V{#�Uҷ�{�}Q���wWձ���
L��:�ν��!;��4&��
C�9��i�n0�����-��٪�*�����w��F�1kz�P�ٜy2�AWZ��A���W�-�S���̰����_)P`��;���E;��"
5`��L�m��ϴ�e��@ڶy�����K4&��	�H�uM��b'&�=�r+�T@D�J_~���4���5Tр��1w��)��~���4���-�	�;��b#�!iB:Q�:�g��߀����!��¾��6S������5p3�ј(c�b�uLS��Us�'�<�����f_��e�<�r��ה��8?���-S4�↹q8�[S�����*� 2����ة�
f<�ʘ�A����[�k�Y:٦)a��M�!H=
��2�ޥ�V��>��������v���C���?�{ֳ� ��7�jƅ��Fi���&���O��8�a�*�ϜS�w��Mz����������t4&��e�+��(�%z�1��I"�Cf�JKg"���P�� �(�j�G�Q������埢D"�Q%[����rml:���E��1����XHe<����:�d���Dd ��2C��^��^
7��x�������M�Ng}����:�]G����W�Q�zϡ��	l�D��Y
�%PrG���=�J&Q�����qcd�ŭ�����2�=~�)���CMn:J���-��hWg������J{���dB�d!D	��5��%S����Y� d@�M��7=UDz$���"32�.������Ssػ{�YRn�сG:�bŁ"�0D�+��fA +��^(�>��y�So��3j�?m�7�M����q����pV�p;�Z���(+:'�J���5�g�n����H��r8���Q]�=����(=�V[
�$,�#0{۞I��8�yt(�nϱ�Z>\�J+*�׍�N�n�g1	���Z���a��7�>t�L�9�t�������5]I�S��Y�<J�� <YP�'K�ib�I��6-�~�c/� �%�.iˢ��w���
^�a<�\BG^ً%�u��|�b<�idݡ.�p���
|�ƪ���7!	Q~�r�qD�}i��A��`#Ŭ��e�S:�w|�
� :�,�b�]�l����؁\Y8�c��᷏M���h���[����6y��m��DF2P�b;�� r\��&�
�k�EԷ�����W�cɉ������)�
��X��%Q�鿈��%�<�}�����rn�7��B��,��7�j���\�W�I^�z{� nw��_�I�c�fv,i�3�j�1�Aʑ��veH��{�0���T�]��j�s�;^S����a�e�S��^��[�lι�"�������#�Qj�m��w�*��%�*� ٲ��3(����"҈ݒ�v������l�k���g!�8}�0��r�<C$����5�{L�L4�����oQ���Jq7iv
�����g(c���U��9��$b�X'��p��M�����B�ء�a��Oŉ����Y/���m����i<�V��t�Kԑ�7ֺ8�*��L-�!ښ^f��A��s�)�9��˕�����r/5ZD�~�GΚ����+(�p)ө��@y���%Q�.d��\�'�Ăsv�z�h���AD&t��Ɠt,���w�m�����������VW4#1��u�$���_Ɠ\�V��i"
=�M��%�Zs~q?����}��P7$�!(�Û'��;4��FMb�t��7���?�S,�:�}�V.�9D�Δ���dh枤�Mg��@c��8^���ՇK��8=��Í ���I�#o�� 0Q��]0��XŴ]:���Ţ����/�z!ܗZc'R,�����ވ�,�M�R���=�h@R���њ޺6Yf����8?5C���r�5��Y,B�U�f㒗�ư��@�D$�tJ���R��w��$�d�����Vd7��ڑX�_���a6��*��.W������y �|�����{��A&ow2?W��,�֭�|?ć�n�r�N?n�"ds���c�@Oғp�ޭ����x:�����{X%j���j9�#_�ͼ�� P*k������D-(���H~܍kL�����֎���̵Ц���>7�!�6|�wX��L��]`�
�D�(��;�&�U������V��a�0��+��l1p^yv�:5�n����7�k�;�!W��p�`D�EĘg��`�5�R���� �7�]J��r���C��f�w{<|�kN},�r61Wb�X����@��c����e��@xIV��Kp%��_&;W�"����!L�怳uZ;N��]��I�A�&v�)�ȴ
�nar�?���'��Y�U, ���`Q׆�(�t	t���]rz�(�n��H���&ע&�������n=�ӝ����Q��C��)��/��8<�.�`+:q�n6��V�мE�>�	&8�?u�^�:��,���L���)Ȩy�?������~ذW�a�t7�}�^$ 35��1�Xӑ�̱��&�p̼jg8��)�$1����<?�c�3ѳ[�%��(q��޸S�����D�W��Q� ��h�]�4F�|'�f_��7+;8�<��y��aQ)B���L{�z�U�c�Gw�$"��mgO��@k��*c���@�)z�Y�ⰟU�Ȼ��5��������V��K~��N���_O�ؖ�z��L�E����
T�S@�	[���[� q�:It	`=�dI�65c��}�3����$Nk���V�4D�V�K��S���!�C2@�>�pۆ�}�Si�7�*���0�a
�VF�rw_H��A��
ߑ98������ϖ'^�K��}�s��[�Ǽ���mݔ��%�N9G�
���xn���[�]lr&�.��6����
�g�������
?ɤkrQAs�ZUb��2T�����!H�Y��jV̽ .�'�n(0vE��m�D�QnQ�T��ܠ��_o�fY'�,��_�֪� .�`58:�t��UɞSi�HT�Yپ��;�XȔ2���m��N�օiԘW��~A5 �Mz"�k�]g#���S�/��C��B46�5�W�^w~&{�܈���T+tF Td�LXQI�FP�)� ���9oޏ��C.���3����GXz�\�<��#C�?�F0*Ǩ��@M!��d��2f�|IʳiB�*��~��(���D�_��dߐg��c�����F��zl1��味��rBY�w�9��M��R4"���	�:Cf��'��ZD��+Vt��j�&�'p
F�2�C�{�F�[FDBͮ_�䓧<oT�����]nM�tO��'Ւq-��lu�Cp��
a���z������ܷo�*��؆0�TaN,�'��&84�糸����|��ƣb�5Ģ�Z<��	J�����9ͷ�}s�X%5t�7�)�(zF=^�r8�Mq2	�`OeW� 3AR��� 9Q"5��hiKb�&��7��^��[����Iڔ1u��f����%��h�G�l�]S0���S��ؙ�B{����5�_3�HIѦ6oc�� $�����Գ�`�8�����+��p�k6�"�m=�ܝ:ڽ&>!�ؑבP�j����Rp��9h��F��@�ڴ�ze\�Q8��$��N�n}0ZE�
Y��������Oc3�,���C�x?���V�X�"���0��ۻ���q&cՕ�1\>.ɫQ5a[�rY����JWi��Z����M \W�{׸��bjD�L�{�z�Au3k�8U� ̂�c�9�Q*�K�.淭P��/�$	ak�#�����P"[#3���9����{~.�
�ik�.��Z)j��3��`�G�	�����Sq���=5����9w�լB��o�ƹCS�T�|`���扭�C֑K�>�X�\�,KJ>4��?�*H՛��(*�e8�??9�.ǅ���#*����,�q=����#X�eX�V٠� ����H?�HA��#��k8�u4dW��r&j=��K_Ef�(C3�#�P�V��N����gm���B�AY.�謒�c�{dO/9G2�h"�qju�&��xO��懧	��@"��ݟ}��k�P����/:<:���AP���O��D�=��1�B;�������3ĊP���F '�-�:r�� @��f�����̯ڽu���=ZV&8��sz�+a 8����/kn�j��8��N�g��P6�O#p����Jp�}��	[$�J��P�i!C�¦��-��kٹ�}#����P���݈�އ�fN��P�4����D��3#x�JL�WU���1&�㿓T6u�
cY}(��7�Ɉշ�s����F���?,K�;A�L&k� mf$#�ɭKVRsd{)�*�j��(�W��,ΤAvp�a��iJ.�(�����f���:Ea��+�GǼǶ@ׅ=i��(�,w`zP�k�y�HM۶ �ևұ��] �z��hY'��2]rLCn���u"��C�$���c�?�-s�$ڡ���;�柦	���JX��s���ٿ
*��~��y�k��GThJpÕ�^�����r�o�������;J�����>ߔ�9H�4C���e�"��ݟE�ݢ����}K��f�\<�\\�29IA��V	v���iO�.T]z<��~Y�-�p���86~&�ɴ:�� �����nc�ĸa<���L�圗 �
�=Ѝ�܋�ک���զ�*L��6��G*T��<�!Ѐ��[�ʌ)(��	�5�_��9�L�k�w�T,��Y��J�)`)[G~��Z��h���ԁ�f�8X��Sd�>�s �:��SK����v�z�b�����
ґ����<ǭ
zܡ<���W'ݩ>B!�0u�-�S9��ֈ�>vX;29řE�5��~�ݫ<���coְ_=+�|y�`@�Y�g�G���:xӐ�H�;2��j�L���'4Z�dfA��շ)?\9�����n��w� �(F����ҭ�A�2��>S��݋�S�y�+2�EA�n����rp�w�|v˺7qazE��;BmJ�;U��Y����`�=�MA�{�ʻI�/�I0��W�X���F�9;�1�	�"�r����]��#X�珇kL��й&��p�q9���L���q�E�2օ�d�L'����.5�m�b� ��ߧ�t�?iUD���ӞÞ� 9�~�l�-�\r���n{��Lh��8�E�[�i?���?��mQ{N��9��3E�)�l~�[�b�:B~k�SFMkؼ'����%��!l�	�E�Z��o������|�y�0-?R�ދhj�[/+���گ��[�0j1)��7���1�@�-����9^��B6b�^�z�����_n�@|��c���#��ws��b��&6WŘ(�$�%y;������%�j��� �Vj�]�������y��\�:�3G�eP4�>F����?��8�F����,3q��I�!��ī8@0T=��{�lA�:�f���\��뮱&�7L�t��E�����߉_��Jmm��|V�NP�{b���Z���}͊����`-8g<�%�E�m��	�h�Ŕ����B��ny�@�3�I>-�fM�t��c�`�޻����j����*�\�{���n0��"�Nܪ4;���A�W�����(��l����:��T�
i�?	���b�-���#��/�������mWM��L�1�|�?�@<�EX��Bmel8?	w��fu�Sfs�<E�Z�^	U�F�37Cӄ�w��`Z���וq��D�(p�[GpS�"Wc��3��0�Ղ�mo�-���N
�zK:�a����ٞ�~�[ɡ����4�e.��x��|Z��;A�ۢm/ȵ����{�'�w�'���P9�&�ʜ�1��SM����S�21{����Q�x�� ����G���
�iP� �@w>��.{�Ӏ�[���\�.�>�9���>Ԩc1I�����lQ�W��]>��)�/�2���ڜˊ�99�7����y�*IИ�x�eYC\�Ѳ��W��m�G]�I�溒� !�`�6L��]^�tR,GY����u��`C�Y��M0���� %^�n �%�Ėl�_�M2٫+S=7++LI�7�<Ww"C]��	�����70��M�ۈ���F��hҪ������?p�� �k-���4|� b�r���Č��0�nz��� Y屰��/�v��7D\��Iu��X���#�Ƈ�:���qW)%�s<��M�澚���6c���\x�|0�n?JI�:qTeP��w��4�)T���R�Qu�����J�}{�9���nH=N侴�@.�1�����ޗ^�?u��p!��I���پw�H$X�;|s)͏P��a\5�_�Pm�_���2 ԩʉ�_=�4Z�9���?�Z���Gs��I~A�&�0ť���2}Љ�)%p��񃯢6��Gr���ә��!��+�]��߰Ӑ��g{�`�5��K3_2?���𜶾}�ec� WKe_������y�����G;c2]�Yn�"�=Dɘj�	IO�\���;���*#��X�p��nN�-���*0ژP�x��@��}�Z�*����J�3/��@�z��
�!��qg/Q�`����-?"�7T{���� �6t�k(�L����|"�669
��5�X\�Wu�@ɤ�c{�����~�1|ȕ\��*|U(A���mb�F1B�8� 	�X�O���� �{�fn���r�Lt�ז��\,A�%�$��{��ʳ=yE�������y5��
�	#s��3��I�4-�\����\� /�XP,"��g�\A�sQ���^�U��"�����\�^r`6}����S�κ0i���4r�{���$�=�(�to{4��zna��{��S`��5'�#��80 �a��zz���j�AS�!��r�APT��^Q��u0}/g���7�����W��#j����5��Rݰ��μ"��^%��o��v�ondp�X�7��9�7>AC��uS�L��2Qn��u-,�H�Q���O���Ԋ6�&0�\}�����LM�Z&h�����K�'�&�ak�9O��udWˌ+T�X5F��R&�:�>�nL�Q�e�l������!v,�~�B�Mv��QG��W��qF�w�~W5�gZ�R�������!C!��^~:��%�P��vsߪb��&]H��xȨB/6�:�p��Ŷw�0�����o�e��3wp�J��u���񈊝U��Y9`�/0��*��V�J%Rᵻܑ:�)�����Bւ�~���̇�6��UEgӬ�5�j�>�\vC��D*.���G����'%U;e(d`D�E��]�a]j��M�
�<��+}%Œƞ����-Ծ�~��x�\���c����us���i��r׈ �����}��hI'l�z&Ho0˸��P~+_��5*"���Ն'���t���뗡�9�Q�������y����x��y��g�ί�z���(
��߉J�*�K�Q��MA��4SW�������*i�)���N���!�QR�,� (� �1$k���i[��7D���yK*�I�>n+׿Ua12;����RV��ǵ[01�ٷ1����67,谡s){�x��/(�R��U���>f��Ƀ�ז� �km��I8�-ª���2x@-��K���9��`B�-M�`J��)f�����R��R!=&��
��[٩޹іo���"c�$��I���H�z��T��^Ѝ�������Tx���t,���"T�=�GBN�<��\�J��)��\۝*�G^{�c���� ���m�[Z;&�2��.�.�9�9XxL�1�����K(+��W�U-��0��	��up�UU\㆞p��ve5�����O�������t+$��V㙋t��B{��7�΅�<dc�7���ZQAj�'8Ε����Dٔ�fumw� դe��u�h����50�����c�k�|��h~�-�`�=z���3?KsW�5�#���pb���K6��P��eFӓ4ߩ��0��e.�1�>�㡿����A$��OtK��s`�c(x����5x�{~�Wԕ�;[���P�d�2��������M�I���V	��Qc�2�q�B�����uhG���ߩX#~Ig\�H����H� S�Ɋ�����3l4��j\Rw]v�%5�G<%y�B<r�d��sI��ĕ�8�_Gv����fd��bJ"�|��� ���<�R!��6�i�u]I��F�K����s�p_�Ɣ]WE=7�=�7;7�:M}&O�f��2�͐������h�A_�g†z�)��os�`���Ǌ1��kV�6~Z^��o��8v}lo�g�4��]ć ���km�����CiWzC�/	���x��nq���gTv���z��`f���*���a3[�z�c���0I� Z^�K�2�
�7 N�;?�T��V\��n2tsc[L_�g�����n`�<�6����6��D�� :�:�8��i�w0�_��\a�c��d���D�S�����։�	��T
t�x�=���P`��Ns���{�ai��n�eC(��L��N��^�Q������e)=lP�Z�^q�O��nV�tmD��E�d��>�5���q1�PɆFdy�s�u�����"��w7�=pJ�G̈�3��O��������>�ޕ�ˆ�URܴT��zۨ���?��\�B��&'Y���Tw?{w��9
=��N���0~n��c�/P�T��7G�l���Ni�$L��1a��0���0Y&��I �4�7F���JiM?�Pڒw�i_rn�z�:����J��Ǯ���nG�9�� R��G)�b�A�[����PO��gh����'�+��a���:My�K�q�����W�s���&�����N-o	�����玣)]V�_�/a{Ύ��[��F'�w��K�i���(�u=/CĲ�����-�����S��<;ѵ�ϻ��Bᒦ��qw0M@
����%y��ٱY�$��"��(5��j�j]u}��Ƀ�4���Ճ���l���݆�q!�Bb��ј�/&�9�;}��z�����}��v�����Z�����<�'�̏ձ�" ȳ���h<�n�K��l��N�N�v��@7)ѿ��l(pEBJ�~O/�k��N9M�:߈C��\�3��φ�E�o�(���+���W8�n+KE5�	S*:�o�7߻~����GD�\�1V��v�<����6@ ����_�W��u��>@[�-{�dP�����u��!Z�V��R�z�7��/P��u[���<������3���^��6��P��uF�:��<XE+Q��t�V}�U�|m�^i�-\�ؠ9�_�k�y2'��mݾ�6��3E��TX�S�m�������gk``1���2^P�Պ}%�}B�J%}�(�� ,�$�S��N-sB�B��ܑ�4	`N�?�G�R����������n.`߾��2�����kĿ��,�;j�i_�A��T�
BA~�}��d�#���^m[)��Ĕ3b �/b�$Z��<�S�tB��w�W��𞖌*0��-(�����Z=C�+���\*Z��u����������%u׶�
����%�Ϊk��Lg���\):W!���,wU���j9�ÆKH��Y��@9}ӧ�u]��E<����/�D��#���8혀` �Cv�b� ����R��c
�p´�8K�����O���1�
QWz.�ɡ�)���y��#�-̉����8���)?�rA/�����0��GrMo6l���2�����Z�M���8�-%����rCpј{��	���=�I���֐AI}��]8�ip�W+��`ۗ1U�����/���8��'��{���u�d�g:"Wv�缜KK���*�Ni� ��3X4�;,Ki�pD[e}��=���tf)r����ec��G���t�JW���� K>�&�D�U�+Q����}#KuO�L$�V��Y��u�
�A{����p�=^(�+�Dma��B��i>;z,��ﻍ�6���$��;�GRy!�Q�(�okU>~J"㜒�3p��GW6�+�tK��+Y�B).�]��s�ŵ�T/�ѐ��y�+EJ���͋��f�cNl��d	ecx�⾍0�O��f��<O% ���:b7����Q1x��NJf�8 ��E)�{q���{9y�7�>
\�R��1�Pƹ��N��ӳ���z\�8��UL�>��´�g�,��M)&رdơJ9�Mv�=XO/O�W�pE(y^�X�j奙�Z�}\����5�0���f+�m>�?̌e�^\\?I��EG�}���$����#@A0[((Tz��������\��=i.A_kҴ���~�k�-1�����0œۆ��7QK�z�Wt+I�2똁}8O�Id�m,��p�g�˾�8��{���َ�Mz����2����
�����e1����i	M_����W.���
u9���X�.1�9:R4"�s`�`{3��A�UZ�A��8�y�������.�1�+\4�r�~Ra�0 ��^��q�Ѳ�i�����є�۱.�a:�՚8_���Cy�`ZSR�{� �@B=5e��+�'9m��cuAm������.�E��GF�����zg�)Z�3Vf�xV�Ak�/�`�e|A�\�#9��+�t;��꽃5�qk��h-r��n�5��Mpc��8 �ٛ�r����BT�}�Sw�j�,�f�[�l����&3��M����O R���=�[)h	�?#��+;��s�5�;e��x/ok���9�U����h��xѨ1ܔ�`��h*�W���F"��"����dp��dĳ���e������/X"vTAY�呖�@5x�<����I���A`�)�<xZ�H;I���l�4T�8��e1�Zo��;�c~��� s�Q뫱Ȟ�5�������UV�8��c ;*����S8G�cS�j�텣��٭�m
�R�.|�{��P�mAD�ʣ:��w3�$n��[b��J��a+�$o_���_�Nt������6�p�����@�M�=P1��c�;���n�P5|��h^�}ӳr�E&W��=;#�"+�Q���Y윒��c��.>�ǽ��'��ULQ�8KֹA��i�5	F�j�D`>Z��<���:x&E��mo�!B�i. !�;���Wnd���z��&��]-�K��1�$�ui��aA�-��_��}ۮ�#:u���!�Q4Θ�IҖ�+�y���O*D�iU+��AT��2
�2 ���+��ι��s.{��R�Μ0�h	b��-�b�jFd��3k�Vv�opҬ����@��ʍ�4��k��E�ł����o�^��MglB	�:g,�!�F&��TB��tE���f�.R���a��<���Z8Mֽ�YxM��>��v�:���B�\ ���=[t ީ�I�(2����۵w�TĪ\s����&P?޹���x�`ށ,^\7����/y{a]Q�Fo�B`�w�1A�G�ͩ@a�e�łd��������
~^d���:B^"��z�C�(�������X�F��t]؝�P	k��o���F*�x�ใ2��?<�h`0Z����a#l	:����y�5�v��a-�����%3E,ټp�7W�K��o?np1׳Q�0a�)�f�L�W����f������#���K}�@���˝��>�7zb?����j��=�-#�])ֆ����Z�x���m��oU��䐿I�,���nJ�%�7����Fk���3+���<�&�ْU��b�NT;+%L���!	�]���Ծ�����0Om�毥�ˬ�c�������:��$�Z7 T�ԙ�EȢ>�p�-I�)��	�[N���m�d����6�b�,%R��A=d���.��RO���O6�vØ���mr5m��"�y2�m$t>��M���?~i@�����K��pb�jf�O���Mg9`f�/�\��O�P���`E�ZR)��G�	�\�pҐ����&�`,���Z����!�3��[:�F�� }u�JIËr35κXȑJ�H$�r�0��gC���>�W�0M���jq~M׼M�k&�<���`�7��ee��x|񮄏�~%�lⶻ�x)�]����<r�F�?��r����Wܱ�����U�|T�J�\G?�v��n���+���~D�����A
8I���h;�:��
2�j8�A��Ѭ����z1����ْU]��+u�DFl�MtӮ���{��?oT���W�z���F�L�z�|�mA����@�5SL�G�9��^��
KtmM���:�\� �m����ɾ �8�o!?29'"�hէG������� Mqf��8{���g���`�]q�A�@���;�^cL�@�>-����خV�Z�Q�:�Ǵ�	��s3m�i��OR��
�?S�����!i�3)��v�]f芴���2���|[��wؖ��v��̽���7���=x��H�U`b��� N��~yӭ&���k�~E��,�O��z��@�Xh�8��~������.主�����۱�_�Df�0jZ�	\�]���1}`=d���?9�f�x�ɣ/�%D�8�d�b�7�����)�Mv��n�D��׊����6!�9�'��}x��	u/�g�������Ff��~�T]���k�C�ԟ�_��)� ]s&N�ڒᛛi��H�z�n �m6��h�VXR��p��y�f/(y�xS��o�=�C�[:��	7cG����d0���"��j�w����1�#��g�ǆMX#M �N�Kle����+~����I��U�� I0�K���>�CW��k�����l�{C�f��F7�p�҅NH �+���$`�#VKͳ��6I[ԣ-\��@r#,�����}�F!���	�l�¨��?���u�LyYL���������j��Š*YD��9/M�`ir<�:7t�P\��`_`�W*.���(};kS":���v�ܺ۹z��`�U��֟ F�ė^j��� ��)��>����aܺ�S����5f�8�B+�tx�7?�����"����T�Y�r/��/L��g��-b(�9�̵��!�>�_Hy��N��2����BK�)�b��>j��c���-*�
t'M�}�;�վWz1�:֥���U~�$613�G���ƀ��R��|1�kj�ꯝW�����O �)���i�rh�u�0����=:����my�
ߡH� ڳ��YZӇ��;���5[�QXV�:�����+��t48�*�1�~AJ�o�N�o���r+K�Ph.�c@�*a^Y��^�r�+L�3�+�Ru��Ǖ� �(>� ���������Mᛂ9���Տ=$t���z�!\�E��vF�����ˎA�����Zy�U4�S�!��#s�R*��Ü�]�I���U�eDo D>_�r��k�O���z�ny��J��Q���ѭ�ӗ`��x7YJ-�tB4��,O�h�����D'[FfNxv`�D��m�?�B����Ȍ 4]і�<��n�_XQl��gaHt�]7�!H���^`�E��nWL"mb�tcWE��z[^�,�X�3�vL.��!�YR�R��t�����C�����Ke�Xp�·��������f�f���K�*�����z�2�v��U*i\�u�tG%`>$!��(#�@����R��eJU/t[�טp~7����U�*@�4�{�E7�-o�����q�Y��u�����{/hN�^4a���橚�3�w1���6*pIdb�t�{����xa�'_��g��� 'G�M�K�ƴZ"��.b�B�n����nJ�vט�&��2�.H2ǿz�îĽ.(����Z���
y\�S�PX{���fњFChm�����O���~��b"�X�9�(��|��)>?�\�x[�CC���jhq�����(>�)�2���e��[W�YK�{[�r`z�I�{�7�d؟�(�����'��0�O��y�8Ŕ���8�U9�t�s�'�� sm�]m{ѯ�8RQ�38����'@��Y"����s�ߟ��p��{�2�x]������qr׳��PT��Z�P���M��9���/�t�6�+Z�Z1��;Z^�?`%^��1�u#����=a�-�X/��@T�EK�qP�}0�4���@���ߜ���:̖�Q�q��^4���lbZp��.�����?;�r
X{.�G�J���nm���	z���M�-,�?ٛ(V'� v=��Zw	~+��*? ����+�C�����)��g6��aB/�O�[,�0��HO ���@���ъcΫ�H�l���祈����'�AVS�����qo3C6�ȃG�P�
���5��ytY��L"D��MĹ� �Xyٻެ�)�팸�c�������נhY�k�[B5�2qS�
��m?ܩ�)̱T�9������U���O"��p(ڜ֖0ƥR=��nʻ2_Bc~)����L�S3�/��V�O����1�'�a��N*���>f^/�s�1�D'�9�W?��ѣjE�rO%��UH>=�k5vp.�%v2n���zI�8���z���N�,�$��_�ۖ��iĮMT���w;D����PM�T7�i�[|O]Jd�+U#om"6�YpDcL~Ahz�9� �MU��j�H.� �b_��F'�cܜ����^8,�qvzK�~S�,S�[;��:���Ln8�T��w\2�lZ0��|�49�%��K{��]`��^j��zɯH�`]lq�S ���ia������߁퀛��#4��� ���|Vaʾ�$ K%��o�&߲�ԣTKVUR�8�cq~�C��^� t�TB�%�0%����'�����6I�b]���ov��Q�S������@��A���X�T-v�*'�޵p�N��p���a���'B&ۦ?� E�+�l(i&�1�C�&�u�@��tc+�W������	�s���}B�A�na2�Jbv
�Fwv|3�����rj2�ĊD���ϝ�����C��� 9�6�أ�ӌxޮ�Y��_{vi�+���R�a��4k����U,ÐNX�E�v]} �r��5�t�x�>�џ�X�u��V-p\�W�)��YQ(������֯�w�H�2�%}ʏ�r{ڗ���	k�D��k�d�V3�1h���*�EYl ��K�0����/�	.f櫧l�Ԁ��-9���!�¹��^KU>�y��W��+E��Mh��_�k�tHL�c3�[���j_
a3Gy���^�x��"�>IǙu���!���A/^Q�4��VK��@tK4�XC���j�lP���v� o�@h�Xv�d���n�T��)W2|U���h7Ah��β����E�UV�::��= yBp�/eM�{�_�ɩ(8�L�\��.=�8�>+�K���TH�����x�pH|ٲ-��o�+��$@O᫮�_m;F�N�rs8/N�0�mI��]�Ħ��ag�2	���*�@��w�����T���Y�9��%=BϬb[r�\
svj���}�#&���`����z�B�vtQ�;f�X�[W�J?��J(cך�4	�3B�<Q�\>��K�y�n�^_��t�m>�8��(��5Ȫ4�#��M��7���5-��#2�Yet��P�}���D'#~���`Et|xkWK�*JR�	-}(��H�ϵu���|�CZ���s�Xr�]b�Ňq( `Q��k���r.o�7�~N�16X�h�jEe�� ����'&�A�����s��]r'�Xgx-�Ċ�}/���q�RJ�#�Y�?)$]��=���+�jA�%�e����O�f-E�%�˓���v�7�j��2��!�j�)s�#_��(� �m��C��Co��N�u؏�9�mC&�ŤD�06�%4�|��hǆ/�p�%��� %�� �>(�������g�~���ɷ��lפ��~�aw6����p�
�qX�~a�΀9���ݸ��{r��N�%�u-�ro�;��7�L5��wހ�*D�����'6w>hp�i�i�C}�;�]�����U�\7���P��uh�&��4��
K�S��Q:c���9��d��%��y������s����L�wn��U�&M�#-,�H�G°w�$����Å]lCz��_�9�#�7Ҁ�栊�Tv������m��᫼���vו�A����a��V��~Ͳ�W�-�|j�(k*L�>��˅]5Yx�J���T��-4@V�u�s���2^��}�l��D�]ͻ���o�h�k�k^h����S��/[G5f����E��H`B��"`�!�_�����}=ѿa"u�1s����	�z�4ZD��q�y����&#���"�U�<�S�ɨRD�
_�wY��B�T {x�5��-������Z�:���417�X��6�2���;��hAJA;<3/I`t�0�r�_�Hi�=�U'���kjW͐�`��>g_a����Ub�I~��k1��UY��˞%� �ն"G���`�.1{np�w"�iG J��?�"r\���4��
�6, k+���ti���b���d< �@��B��ҝ{ P�O��Ez�b�+�!Pw�#��� S��S#E�iL�޶��T��~�&�ho���f8(p��?qS�8�aň��@�-�yn�.ݴ�Y�Xp�Dی/ЖgWV����
��h+������@B�j''E�R
4���%/��o}�ɀ�䭰��`�1߫k��z��dO=��y�D�c���5)9�MZ���ڞv٩�DԈ�3]ؓ1_����yj��!��2�2*�V{vD��c��wT)���Qq�PD6䴓�4�s�.8H̳�bMz0n\I	����
Y$�[zG��A%7G���z�9_��p�G�����X�e,	��ٝ���=��1���>�}/�s�Z�;A-��n+�a�e�v$^����	0@y-�E�$�nT0U��p��B�v$?��͵Lo竇K_��j�>���FD��#RM'�p����TmN�yL �lyG�fsԬUZ7�~�q��K���]���
Ah[Z���Ʌ��r� |��#�M�entÓ�XY��<g�3�ݜ�g��.|^<\��[{0�]�h)�r���g7Զ���%�P�&�fS��|��>^,�hH��~�9>�FR0����`�T���L�f�����T�I�<�3V�*[q ��a*��5�e`>���+�$f����9eF2Bi���1����I��&��`� �O��t��k�;D�Y�Ui�#~�\\5T�X�a�F�e����_;�X$��Sj�Ȫ1�A�V�����"��)v��M���.�;�(t�/����8�{ �;^#Ó�evǸّL�L�ϻnD���up���V�~u���
��{u����fm$5Qq6{�wm��Չ{ � B�R[��Bz�c,���LwH��8�2^�N�� eF:�pcP��y��J`h_�T@t����M�Ac� �-3MӨ��,�X��pbŮ2��'�����ƢX�_���j�Z}���2?J!=^<�6�w�wE��H3�9�	m �p=����3��3�25;8��A���AK��( :�P\���qA�%%3��zt�*2�⑞�����+,��b��Ic��QֽПmp�s���C�Ov��*��38yDyBɶ�l;��u������#��{)�� ��r�<$��l�&r�J�D��|j�><����ql��2Sf3�J�����8�E>�:V����h>g�m�$��0
�|����|c5��OABywG�ʧG�����@p��(�8�%ǔjC(�%�5��CA���yR�KǱ }�l��On���<�h�oO�p֤����l�`y�y��ƶpmy�jK6��a:�)��JY�X"�o;�� ����*�_}�]Q �4�ᤆZ<a\���(TC>�T��ر	~�l�D� }+���	\@T"c��b#}V��A*�m���Δ�3߽H�뇴PIz ����]�rc�Q��ʑo����C�8������H��o��|`IP!�Ҝ��H�@�l� ����#�����y�^�ό][<m�(�3u�Tp�������>Z�v���O�[C冀���M)"o�InZ�oT��"�����	��kX�^�a���a����V�\����a#�x���0.I��~���"q�ʃ.6`����wa���.���1	�g�����KW�r���/f|�;�^U��Oٖ��!�Q�α��í�(�jϧ��i���LD��s�f�+��*>�@ �Ӭ.%����������?�Dr��&'~qKs�i��Ӆ�I��"]����R���P�GDV��PclUL�תgA��7������V,��1MC�;8���]:z˕#_*�*{�@P����֠�Y6[K�1 ��5�s���TR@��� ��滍�b춵q�p;Cj��� 3�ȧ��>�d��DQ| �Pd�h�ݞ8����_�%>e��ᝬ|亝[�ޔe�o����� ����fb�ɩ���W�/ӪÖU�1�a���Y�������O� 6�xh�*�r[Ϋ������Y���".ƥ*��/�*k(���xK鈟�6����D��I1؁1oD��ˆr���ҽF��;F+ڈ�1-�7�qUn����!�m��JR�����<�e J�I��\X<��j�%��w�um)�c��bN^��n*9��n��A��ZW��mz
K�e��Fו��dt
����4��pM�qw��b���.o�����A�~��*nhh%g3l��xZ�W��p1)XVA�Zx��ٱ��pZQ\��;������L .�KgSz��
��K3>�UӴ�����Jݸ+31�h��K`;ԏ��mҽ趃/����x��&z����9k�L;KP���}خgKd{�Xx{�r����m���z_nr��a��0d	�^af�̧�c�S|�#����}�0�<�L��V_��i���y�w��H���� םv�9YN�� �(����%ǶE�3��3�aP�X�֦`B�2���w��2�{E�����"FwY�M�#
���t�r����G}�oT.	�-뀯�Z��`<�v�YKMy8̶�̋sM�U96��RȧC���)W��m�6�14��ß$�F��� ��¹v���Z��A�V���]�o�J��T]���O�S�����1P���e�Ϻ�1f�XwE���GXn�f���d�M�.*{�]gV�1Ki��.lJ�2Oj$��ro����`�;py!J�k�i���A]i�23z 8����Ͳ��q�X�Ts�;5�� �)w����m!B���Ƌ�	����L�nb|�s�t��U�2��P|i���W����}F�:o�?xa�+#AF�،��4�ǄK�j	-J��	(�Ȯ�Wog䔐v�ݫ��=��M�ږ=+�,nY��\� ��v��Y��A�bj�7���f�HE��w ]�l�"�GB /O�V�]���&�W6�e�O2W�,���=�8����ZkNQ�w���9�*���A��HyF��<})&�Q4�$��pn��e������Jl�3�6�^��~n��~��)��Ueۡs�7V�U ��cGQq��$���i8��E*W���� ����w���A��1c��Uy�Պw9��jr2=(8�,�O�W�J#q� �X�Ȏ�ej&�*+C,����� Q<tُ۔�xq�4�n=����V�#&a*Y`# �s[�F'�Ӄe|�6���G5c=Ycm���kVSȻ&�E���3���7<�u�`kd:��u���:p��g�ӫ���G}���f�*S���M�������& \�$�Nd0m��O�^�O�*�^&	�x�We��H�[����{A����޿�dU��n������K�.ؤ/�i�{�Ƀ���I�dir����eu�P����sh��.ܑ���}�DE�㚇2q!�%�Q��h���|�(�'%c�s���D��6�g�VbԾ�R��9C��p�[S��:�h�ƍ��m�:۷p��F1zhN�{B8\9��l�dy�DY�QF2@�W������G�e�{9��^k�����3z�ϯ�E�̨$���t�M�q_�uj�V^���Oq�(ߥꡬL�������߯u����eDnl­�7V��y� ����
ػU���RA1T�y���s�)����"�*`n���|ET�Gߛ;«qa�d�����S�es�r���j�Ah�\ҽ1Z!������5��$�G��	t�ح"�4�֙�lM�+Fm�Pd[�,b��3�c�G"�?(�n�J8[x�.�{ ��<�B�ȅȢ�\$&��������ߜ$qW.�zV�|�&$�{�K��O�
G�����Cc���+T�MŽ4����\ N�!�7HS�j�"ۏ�'"C�V>�B�����{�'O������w�,8�F���]�U�����N�P��������=��h+�0�4��y��o���O���q������a	%Q���r�u"ٶJ��m������Hh�� 9ĭ+o�����B�����o����$�|I����~pa�>��L���g��D7Op�h�hA��U�"(.�^��*@ٶ����7�$+���M�=x��Չ�٤��n\!D�?6�3Z(L�Z�S�|���98%�64N���j�J�dq�z��fZM���®�2���BĻr��[�d���GSv�Ϩ)!��>?��΅B���r��Mr��o��Wb��0M�JG�g��^:����*��1�����.V�������gpد�j�:{��R���n��h^����y��=-om|�\�6ȡ>�so������R~�@�J���d��X��H��u���S�ü�,ƚ���^�c���$�����t-gLNֆy�j_�u�RC�%,��䟒q���C�!]߱6PAb��翮�w"���:��*��f��#9��	_�_ȁ�S�i�2Z��59I���YYSM�������K#V_�{�E2��zA���Ϛd��T�$)Ɩ�U[�N�Q�+�ϒ�QI�O�׈$>8]�!�a�0�+4�q�L�.<�E��g��;b�۷}9�P?��gs�.�'�Ѧ�ғ���}�ty�_A�Ar� ��C!.�OS��?��U��P��f �n�#��p��=KUX�^��I*�a� ��i��~���1�-Hh���2�v#H�La�_h��"q�}�Leⶅ�1��,VPT"��r�f b�L��O/o#U6�5��w�ޒ�5��c���=��k��獉a��D����hn��pA�O�n5G��<,�B�s5���P# �К��q�����?�����3��D:'��S/c����Μ�
���x��pai�,ES����J��L���V}��E�����}�U�T�(�m��f?e���u䵈Ru�֗�7V4����M&S�]�߼,��=����m��C]R}ˢ��J"ӳ������H�K#����:�L�e���]P�����N����$�o䓫3%{L���R ��0R���忩@/;d�sp���{�A n0��"Sn�*���Ke�0r�����O�=m�mC>Q��t�)�_��n*^Z��xI4�(�ur�ʓ�\��+Mқ4Lb9�a�؜T�����&�Z/����r<a4d�z;�>�o$�o}��O�I	�}o�����U}��[E�n%��!/@���iz)��|QW����-=$�u�e��m�'	P�d�g
��|'�cw��5�>5�-!��E:ʊ��g���T�,��A+��;#��V�9�5j��䶩��@�>7��\6��L	��V�Ց��Z��8�£�O4@��	6o�+�QB�S�s��ٓs7̋$n���7��;�&~92�H�&P�LX�A�g�@j��=ަ�9▅�M��k*�2$�R�ӯ�b�瀬�A��\��(��S�o^�������׹���"y�WJ�t�y������qإ�(܆�e4(h��W�A���7�G���*_,.U$q�� D �59'N7�K�ZU���}��XG�7
k-a�me�]���hQSxUr��9[�c��*30�j��^��f�[��Gq1���0�J�S�y��㰛 @:*�E'赵�N��\���N,���1�\C��q��6�:-�B~��04����P�F��"��4�	��~��,�U��js>A	��0�E�R�|�|�𢶸=!&�"D"�",d���
<�t�҆꫇q�l�rTڜa�-_�������4���1�m�a.�Ɖ�jT�0�m*B��v��!~�Y��:�@�$9f\�rN��w��g5n�c���"g>���!�G���2��?z�_s���&��������NI'M��K�+[��(��O�1C��(f����E��� �L�R�j)�Gy��I��Ӧ<E��ܭ��7P
zުy�W!R<�?ۘ����[
;�,���!P���Xв���hPF�D�Q����\����	:�q��g��$}c����ŰQ#�V�RG�E�O������R@ a�a��d�c�B�
f���3�N3�s�{���A+p6SaG��&څ�"�������{��Ku�:j9���R}Ne����lg�6�m�vZZ���&W����8B�߅�L�xӡ�?�>��=]k>�pZ�yN 2�,f'����K$�ZNO^��҅��6hk��|��c�IvZ\�{� \��?V#�g%ij���s��.ڜ\�le��s��	j��1K�ܸ��'�.(�f�ym���p��
S�>��A�[�Z�|��ݽ�/����쐸��S��~�m��G��Z����43�id�)5vT�@]1��"[����t[�'��u3I$¹5���pL'T��F��%��A���� �q��s����|�k3}EлӪ->����t-l�7�a�V�[�'�H6��T�%�����|f���U�X\�n�!Qޡ"���� ���s����+��ۼ/uބGn98F^�fe�k�:Ft��F� $i�������xr���KӖ����)��9��f��'_�a�K�'�]v,v[�G��ڜ�LKO/��Z��)�w��򐼑裺�^a�{�r��>�v0�ё^_g5W<Z�6���a�1tV�W��dY�|�(�K'��z���]���$b��n���A�Jqۚ��otI�d�G�%U�lG��3G�W�+-u��d���F�գ�x0�<�L{�l��,�nY��VsC:p���K�' Ca� �o�l�K-�m[�(��1y��s��#��+�`�N�)��LV�E>9i)�"��§J�/y�k����U�l/F]̯�@����o�81sѦ)����]ڦ,y?��OMΥ�;�9ޅ����M��z���F�~u��S����ˑ}M�1�byz�,��v9Ķ��x[��y[<��ж���`2�I�[p�Bh��\3���Den��[��DW�]�F����ӥF��W�/�š�g�⤇Z��}��T��Y:���dj�6;w�RI.Ny s�~��-���MR��C�G%.��2H���6#>����U���3�*�l�DCd���Y�dH^��B���qC�e,���u�!*8��Ӎt��eH�CG��ȘvA�@�}� c;ތV���]�4P%YH���,�ʤ��ð66�h_s����҃:��@������z*���cQ����X��C�����@mϗg�%͔�r��g5)�-@S{��'��;4(F�o8N���A������K?p8C���'�n5RH��[\��Eq?exҏMԙ��@v-!F���`�]"ƕ���������^Bp�F�;�&�.�����.+s?��ţ�6޷{7��6�y[|��<Y|�V�X2�����HسbDCꙓ>�!O�����?��/��l���C$�d�����.2��Ȕ:����1�ؐuV�2{��U}%���E=r���.���4��NG)��Va]G)��<`G��1��_����ᶕ0�]޲�|����3������˭sJ��&�WD)�^@{f�-��M�^	8;�|�~g���v)�q3H��AL܌QbZ�vנSHS��}?�)u�sy�T�o{:�l�
s�=J`{���r�k[�T��<<���>uu��OQ4A�GY���I:_���7喝��w?,P���W �A���9�a��%r���U�d���g=Ԩ�;y�u���т���%�??t����K��6g9`ޫ�X�a�>�'�5Y��`�OM�t�oZ���S8��t"nDp-�^��� -0�iH؄�[�y̌z�&��I�jml����b,/B��ϼ��G,R�A<�]��������%�JL���PQ���k�yE��dO;�Oi1Ζ�G���+,4�C��P_(v�E����L�G�`|�E_D��7txL3"j�xEU�7��D����ve�����0��e��� ;2�kpe��y��N7H~��� "Kp���J�vLd17���61�Zi"��!;e9�	��3��P�8aALFz�4C�����~Fߋ���%^�ޞI��Z����M�ڒ/	�eA�6�1g.��
dv0WId�I�Wo@��8����t3��7�j��W�� ,?����h.�����|�+����n����v[S�}�'��8��l�J�x���:�f/,N���0mH�4�� ���J���N�n�E��@�WA>%,d�ku����C������ryg)B�������Rj�+c{1"��{�;�1�i*ʔ��"�a})�%�E�����,'�}f|��@�ߚ�ś�"Χ���I	�%��o���O��{`�x@�5k'RS`�)ڮU�Ó��D,ɼ{���M.���E��r0U|�'���~�_�:l'�'��؋X��R~c]?XK���wgn�!�{h�q�n,B�	'�5�o�S��( svT��s�̎RTgb�@o4�g@P�c�o���Ck��v�'VV�B���s��d��)?#��p+��M)������wO6��9��Z�%����g�\g)�۬
ӏ�T�:���v�)t���>��%��f~�:���i�i��miS��B~Ĕr�c����CF�^�ԁ-��������q�=p�R��yeΘ�^%�阮*P|��#��3~T��6���� i�{�o�d�(sޚd��L���ML��;��ἄt����h�.8w�� 7��?�u�m��U�SN��擑��ݏڙ�:p����H�_)�Y�W�1�������lF�����撴��E���B5˹#J�g�~���Ӝ�t�Yg-��He�tk�R��,{��-�v���\g��Æ�8�ݪ�9�� ���ۇ�a�� �hkē;�������8+�r)�5)�H���rI��fHo���)Z��-��S�2��qs�膳_�c��:>�>d\`|�s��!=��n�:��9�38�`w�E���`��{b��Vv�ߏ�0ym��K���h�Z�z��Q�C73]p��3���ȳv|4�E�J�t��w�ms�[��Á�e�8;��@q7/E�U�M�鍽���F�᭹?�F}�&�ӗ:�����-k
��WI�$�aM���(g7خr���9�G�H^����Wi�Q����)vFuV�$=�]�1���eu! 
���x�ti��/0*����~�Ie5��oAr�.Ce5��hzw�on?$<�[�`eUM���� Ďo\���,i~z�����~����h�b��V$�(�F�$ә� ���0�}���"���lJ�i��z��Ǵ�0�DF��]^m��V[��?��	�H�V�c����zl[~מ��U�1��m �������e�ll��z\�%bH���!�m���,Gu+�����گ�3�`Snc<�~9J���|W��-&�x��K�r~��k�YH�^$k��7�U�v�Z��>z���Ӈ���h���>���`�H���IVH���X��'�<ԗ)!����`^��$K����#��zY��n���P��ȋ��5�Wt���h3vv�� kĩ�Bl!�~څÙ��i�1ݿtS蔸;�l)�[��Rpo�������Վ�s{���(���c68�:3[d3J���8$y�r�|�!�b���_~����*�U������\K�2�Ԇ߷Z��|ݽ�
>ν+d�����v�&u�����EH���4����q�q�����6�D�|��R�	$:	�P�Li ���V�;��iw�����Z�����靣���Y�|��C�Ҁ�3�RAG���!�U�m!��V$� M��j#b�����
��0$�×V"
l�g}��- �/��(�BQJR��5��Pa�E@��=rl��c2��}M%����&��~"��uW?��}:��4p{E�i����y��Ҳ��_�$���/c�-(9���r�Nd���2�G2�V���̟�r�x{}U�r��ŠN��k6��'�$�/Õ����{u�83��p�۴i� �7�gf@������RL�
��@U,0�,j���awW�m&$+�ا���d��z�Vg�:��&o@�EUw�0z�L4�워i�b�֦v��=�fFۄ�X���<Xj�PӚ��D��`x$���sX����d�ʈ�{4��@Z���xy�K$O� Ӎ���`U}����0�4����r[G��DJ^�[4ݔL�������6�Q;�%XE?K�
�q���\�����x��c�t#��5�/������(�?r	|���	��_���. �o �C��h;��%��}�t��[�g���i"�����T6�M#"�So�@ ��7tr#O��1� �?\��hs�ch�[����!��g�XoU ��^��GB�e���ߨ���|���o*�[/�J��C�� ދTl����Z�ƣ;����z[O�_u��-��BB�XB��i�<'�yoP[���"�W��� �s��WX1� �@F����tb��1v!� ��d,n���!�u���+h�T�4��w��Վ�������܀��¥R�{�1��|��a���0�-o�=��$�%ܖO5���=w�V�-�!f��q"&w�u҇��b��2���!��/uEy���LD��܌��:��Gw�[�u�����?~�V��)�w�z={���z%`G�am|�{�t�6�"�af������ ,;���1��
�6~����Ե�m�]�3�2Ů����E70��*��\z{�I�71�"�����:������de�󌍌'C������F� )�dA�g.:�-1*�B -���cFT$�9��@�;�4�U�>�S�ސ��Ȼ23�3�sk�$EeזF :
V�H��cj.��T4:QO��@�����ǧ�q��L�g��WM 5���q$��l�Rtـ����4���� ����N��X��!>�gYr�ǣQl�z�R�����!�E��uog�zѴ�����!�A�QH�(+��Z�HQ����XN5���$����BT!�TT�:&G�������_ݑx?Ї
���������]�=G.-�A��db�Zչ�R嬙6�뛯uxˉ�����\���z����v�t���U�YN���Mޡ%�f��щd�w���f�)�a�`��;��i!�y�d5����1 /{��z ��O��#�޼#�A�������A�^�]/��jFC�进(�2.J��i�ŔhŮ:4�@'yQ$� �cQ%�c���{�@R(�#�sؑ\إ$c������(3`w
��:��Xzw�6�B�i� 4�]����9X��@�?jݥ�ws�/�,t��r�q �P�cC�YNJ��U�������f���o0��$��_�j=�هEg�H)6�����m�U�:��R����?�����C'�?W6����/FT%���op]:0����GC$Z\�K�����`%��"�i)U뒖�'�X�{���3ZbSi��%��ʚ<t��P�`��& ��yL.�`哂�����&T��_�ܘ�$��D^ĵ q��G)̥`����`]j��~��l*���`G�iMlo�Rs�K�uB|���ĐUq�׊�H���{
�a&�;�3�6S��o_���|����������Ԅ&�H��8��<�AAY'�.l�ٔx�؉��:^$��)���@36 ���C�Z�&�Z;�"�.Ci[t�D��p�q��7�+'GL�r���w�5���58
� ��[�����-��&�62ih���%�c����[�%$B I��R���ю�a�;�n\{֘49L!�?����G*ro��S�C*���&8����Y�,Y}�<A����T�T�ݵ��Yq*M9L�=Z�S�D�c��c�=��4t?YGĸ�SLp�w��⤑��\������zQN�Z�������7n����n����=	�S[� �� apII3t�lgL���,M��A�mIpȥo�AvV)��"�4�n���_l�h�X�B*t���\�Ϻ��n�z�0*��,�B]9D7y��9�3'��UI�-'��kr؅U�Qj{�{���~J𘱳�S�.�A9x�,�*tN����8��u�)Q>7	�Y_??�@���j�U�|m�%���@|*?]�Y�	������)?Hus,�*�ܶ�����k|������s�T���Ex�F�M��h�p^��JR��6�`f�مƜz"��_�WJ�G�],l�u���xaJާ��pja:�?��%���p�����Đ���ŉ1.]���c�bZ�
�[�ÃL�O�s&�&��Fi�6NnU�Jw���_����EQ���\���0	�B��2eV�b��o�~��!i�ѮS�7K� �a�3Ů�����0�xw|��/�������3| ,�a�Ŋ���8d��P���J�:�L��8W�a�S)�
��2]!�K���.@����q�
a��e�I_E��s�ә�ܰ��0׋���G��W�Ռ��U��3�e���H.4b6��Bh�`!S����-_.i&��mߏ�!�~��"�s�*N&sϞ7��-��
� !�g�1�t�������@\{�
�ߜ��ѿ%*�����&/���-�}�����!�D��I��'�Joz̡�,��$���\[��;i�|ы|�la]dv���?@N�E�x��}&����A�=j�
�\�����qw�.��+~
�E�>��.����?`>��0B��y�{�͚+Fo�e��,ay�#������sz�ן��`��{2���ʡ?A�SX���ń�0 ���XQoI4�>����tU��W�Z�@���Q鍊	N��o�����#m�U����hܗ��>�~�Ϭ�]���t���R�����2�
����1L�|���2{������p��^T�T�4/ŠG�KJ{u�rLN2�_��*�ӤG�el��M�E�+���`A8�yX)6���hp�s�4�m�Ns?���������Vs��D~�}�4xc�iRJu�G��p ��b)c�Y�JZ޺&��^�Hvm�kE�17�i�����4��L�d����� A�;�t�!���Y�g��n�bdc�okX�@�1�Ǉ�h�r�}\u�x�=#쭟/#Oaf�������i�L��m��Fh�o�P���L�HY�k�X�Zf�a�{�E�7����W�[����@|&!50Tw�QC���tɻyU�r�%�Lⱃ-m�K7U���(�m��∋��X��Z��TΗ��=D�ؠN�D��e+ v�P��������+pj�u  "�UW� �����OZ5���v2�VZVH��9ΓC�2�ޕ�߬X��#l'p�A����~����2(�G>Ԛ�M�!zt��*�C�j��G_v�o��3���K^�L_�]��R�sN�!m#������p�� �t�����-�.����`4
��,�;c���&�Lڗ��J�Ի�&�p,����s��9�^a�v0Ui�cXy��Q�t�.!?n& �Č@�T�HX��r[�mtл��l�^�kb�s�C�К��2��p~c��|-�����GO*ou@le�3B�E�x�(��y�I�P��+�;�1�XF�R
q$�P��h���9�>���ԝ�b���@����6��f����)/�e�8 }���%�����%�~0笎�b�������Ύ� ��(q�=� 1����|J4;�3��if�0����7�w�#��޽]�`zB&�7�,���6vMI���5L �� ��M�H�x���{��h��q�|����2A�#�#%�q������8�yc��I�H���hጿ9�[�G%uq���A����wd�Xgj������i��t�X�`���QFRi��ߩ��:��?�, ��i��`6$ōA`�o�\�D��FQp��G������X��s��G%���\0�
�ɷ��d�2߿%hۗ�JQ�pj��e�C���t�>�s9ͺ4Me�&"U�
_�:�py�6�T�HAjڍM��zbNG�p�S#��s�(�S�N�8%���74�0�4q���I�C>\����䷇���PVM@��bqyu�6&H��)�ӈ����+�����C̭�������"����A��W
t+����e�+"�dƮ�aҬ2�L��5��{	�y����������,��8g6���b�U�=��N��雟�)���l�Luq�#Img������VGZ<�}�a�o�f�3��W�C��n�.A�r���&'���^�*(��%����dA}nٸK��eg�w�������i��q�%���-V\�ߠqZJ�,���q�Q]����0"��3�2=U�S�䟆sO�r�]�8��MƂ��+Nהx��"�o�N�|Z�q�3�.�=D�k �y��Ί9�set��u*%C�	�#w�@�n�@�̂P��[��$6��p���ioL.>ˆwl^u� #*蒃Ȼ�y�:�鐤ɐ���Zpq%x�����P��-�S��=j�k��z�������n7�w2}Q[��_�V=��t��@t:��3���dt�&A`�R�e�t�oȪ�3ӝ��#��x0勚���=P��t�;]�)���gz���#1�����7��_�
Ar���ߺCM��֏6Z�@Kc(o�s�U�'U�]q&N�׾����C�%ëd�ré��rUl)�Hx�� J�U��0��D% �u��r�9[आ�غ4D��;��	,)��U�~����	�s��=�F3yZxS��m�I��ShPQ�֪�_��p	2��#�Rc�9�V�!~ͽ#Hj�ٖ���'�v2�UXu��G�E��Yd�u��Y�Bd

�g�<�H)�3Ԛ�1~�N	P����)�X���9��Ֆe�2��lIYF�2��pI��Q6�%n��Y�O��%ߜ���M��1�Rn!���{���9l.������{�hQ�T"/6!N�L(�K	��D�&+���8H>��*k-� �s�$O������an��:[~e���Z����Q�8@��=�p����
⟆��u�#
9H�,�kZ@���Á�?}��<y(�J�1oX��͘�M6�N!6b��#����T��v	�dB�!1��x�}Ċ��wA�������(���ۆ�(y�&���p����l�	Yo��yk��RJg���$3L�6��(�Px������s��ݽ��Jc�b'W@���ad=��fw��)��T۸��Q�I���2F�,��k� ��'��,�tA�[B��uE� lk�#�cn�H���ͤ�*�'�_��p�3Z57BE<�Oѭ-� �B<�p�λfq�\����c��D��!(-��BA���[TJ=��+
�p�VP��`Ȝ14�[0 <']��+�3ڂ.��c�{�t�Wb$�M	bh�Q<��ZGq{B�� y�,<��S��|��:w��Ø�T���ű
�& B��ĸ`5�����6������J		%g����ɹ�)t�'�%�L�;���p�6�YO���j
ٮ���R"Λ�>|��dm$}���~���Q�����|���6b	%�9��<���d��Kd�
鲥���ܐ�+�9����ڮ����I'�̀��oNe�N�amcXs`�����x�в}_�
g͖������tJ2;ހ\y,K�z������X333-;�K��ڋ��"��e��Q6�"���'N�'���)��ABr�_�a��،�S%�:��o٪h��L���)Vk�U��,�f��C\�6
�I�~��"����<i����%q6���u��|�<a��fذ��!8Sˆ�O�i/�t[�tW���qNo��!�3%"�:˩({�ruKx��3�.��L�����H`����ݕY��<����J=�`:W��h��6t����6�������_G���pV���j�`/lt����f�5V� ��l'�vE`cC�Q[X�hf�yn�>��li	�P�1�-���j�e��P���p9���͎����nCCY����˸h��;��c:�ϔ�ʦ{�&>R��c.57���M�|��u�u��Yr�gL�hj�R�B�/IK�瞴U��{����$K@��vԥ����B��������1�J �4u�Dce8�1l��4Y>5-��MEt��xb�\������zj_g`�[�`Ղ�?�#a��J���R��pr�0��q��ܛ���-�_n\RWEӛڏ�؎b����O,:������4S� �^i����C�r�vd%�"1�T�i�TJ2ɝ��W;L�mq�ua�O�Ta$Ϙ �m���)��2���)�78,�P�{��~\��ʎ�K��=�AF��CX6�W�y�-� 
i���9Φ�4�b���w�N������}��6�� ��R|�Hb${Z�ܬ"�{��zO��)\�rmp��)Yv�6�N��&���l�����JiL
�QßY=|ٌ:���0��_q|��h/�=��2�:�\�?��g�,��*�[E
��X���T)�斺�o�Ӊ\�\��HO-��i·�{&�ѳ)�R|�-�G��"NN����`�$ �O��l ��1�¨Z��Y���k	:9,S�EC���]ж��|�!q�\v0c>9�{���M��6>2`��2�+��q���������x��K��〴��]<�vX�t���X���r�Z���K�9Ŧ�zF���F[&{����g���m0�R����l��#I!`B�����Hե�Zрw�F�T�Ot;���� ףj�X0Z<�o$!y!;��\Yu�ȁ� ���L㺂�o�ȑr�1;'�P�2����+Η8�����WSN��5��H9D����b�%; T4����}���Q�f]����/��[�"����zKY�(��\oRR��F98~��5y��ʝ<�q}��
	�]x�k xy=������7�4Ć���r:qCIS�Zz�_�)���v�sB7;�, ���"A��ф�����!������8��r������Piqlܛ�d�υ����E?����|�)L�4}�C�Y��Yv�
��^
�~��a��F��e�~�x��fnKZ�r��w�j�/)����4_~����_��r~e�!�plvE��v��K	���<�a^+����<�Y���e�����j�J59�
��ʱ�eҭ�.��]B7�z�X5�f�,��_�����x�w� �G��Ix�=���z��F�~}�f���>��@�.�U�l�|��ǂf#��Z7��n����:c�Gh��j��Ӌ�'lP�u��p�]���_��r��tԿ�����V� ���@���:��e'6��+��dT@����%Ѳ>XJ	;y՜�!�Vk9��!\й� H���o��mcgc�����>D����o_.�����I��`J̜�Q��#��r�b��g̃�4���plF���Z���J*�q83|�?G/�4{H���^4���sOS"	E-��^���M��˃c�NR� �\������:�E!ؐ���u��sͬ6Ɖ� .��3F�2�.����[�v�*UH^�bO[���60��_��8�w�-~&�ۇ�w"��xA��N9-K�#�����K��
5��������y�6�Q�|��Q�e㿆<\#�09K����'6HU��؊uc۝����ݚ5�� ~���B�~OW��GTH�*��&Ȱ�8Ǟ���%6��Ψ�nA��,(��֢�X<e<�݊�������>y�����z>F����=ɵ�w��s�{i*s�qh����Q�����ᖄD��v�%���$g�j��h�O���N�~��Zi���3�:p���RS =[��f�p�̨-���IwE�K�bE�l��1O�O?Įa����r*k�]�����VGu`�J����_Z0���-�M@t+��g��O���?QA��ߟ������Q����VI�	�n���$�����v=m]���:����@�1��������L4���q.��Ŕ�
L��5�/&�o�z�Jb�U���ւ��MS�,������E�N�^R�e�y��}��k��ζq����͒J��+G�Ѯ�1�\�e�*��Tw�;�(qsº!����++6ݽ��5��{����7���.�L�(��Ǘ���7��1txXX����!���G�^w�2�փj��)д��t��M�Ns���*��e���ˑ�̚�c�^`�5��U����/���B�x�Ť��O	�C�R�Ҁ$"EzO�&��oaC׊#�ISiw�}�r`�u�Ѳ�|��R����$p�߇�	�m���x�B�q��*hzC��pp�o�=�w� ]�
��.����7?j�Ȁ�+�������� ��"Q7Q�A�#�Ì(�e�
?BadU��ɟ1���ʄ��Z�4�r����51��sz��6.�3H��)i�W'��8wƿ �*jg=a,%��9��4�-MX�xR��
A�U�WF��р�=C���)-K��1�e$"Ŏ!�s��� ��\=����W�1:o{�8]��7�C<K�eV��8�o'?vĿ8����6��p2�&�C�$&U�FA��/�ú,�"1��D&`��U%����D��2�W��L����2N8Nk�������)P~��65���[�'#ЉZ�6Zţ�1�	d�4yx�.�= 3�6��X^��������>ڢ��mC<^k��!po�\L�o 2�kW�D����ln��Ϸ_J�}�V6�R��<�+�&�iC�޷��g�I-F�W>�zÅ�"�W	;�/MC/%��!�0��f����\p���r�+�%�|��S�4eY(IRd�� �l$ޫ��v���0�^�v�Ⱦ貌���;6X�F.�C���*/�c⟩[$� C�:�<�����1n4_w�7Z�D����ͺ٤l�㕌�|a6lT-t�F��/���Vѳ��j?��ܟ��Ԍ�Ai�Q�=V�0Nے�Hi��˰R6�s�:�����n�)֯��?��>����}�	ϻ��a<H�������	�=��6��c@x�?/>v��>����2J��uv-����������Y�g7�.(��3�=�^�KBR7��<p����FiHة&�����Ι7V��'�at[��|���� �::�uC� gq&�D���O��cz��Ҭ܋x�ԉzG�!�MK�i� �#�m�ń_đx][j����-���z8�m��Ж*�1�m}֨
�	Xa����>F*l���{\��$�t��ʺ�� ��x~l�WBud׉�?�4������vhq�	�k�a,�M�n��b�Rj���_I�L��=�� ���8�BNt�8ݫx�=��q��;ǖI�@�AVX�$?�Ȇ�u��ݖD߹L'k	���ϗ|��跗�%]^M/�Oy����ܧN%J��Ļ#[����X�āZ�pP|ٻ_�@Ɠ@J�,�t��cS�ȥ�Pi���R1<j�޶1�	`]u&�Mu������I�;�S���� K!��¥l*|:Q쬿��J�ݔ⛨�3*��7��K�t$~ڈ��M��*�b��䒚���ZA�J~��+#cJ��Jk����KC���J��O��f_�����8�q-�u((j��[ɍ*5+��S[�:��ڳ��@�e	��P�����}#N|)p}{6\j>��e	Ӗ�'FKs�g��[VM��!��E�z��re�öU�@��m�()6#�s�#��ߠx1���R�#/����'���JP�/mp���J��D~�+<-s%��� n샙Q��[D�)��c�=��
��Jd�0����pg����Zyk���:���i���m�&{���>WY%�V��ūT��}�������4�L ��c%[8J	�=�F��6��6��4����k��^S�vI�m�*0�w�����yOV+�ֿ�w��/����N����E�k�1����>b��(ֆ�CQqo�!�b$z�NF�����	Q��'�)W�c8{M�tτ��~��w�W�r�'���wv{+N��|��?$6�eh��ܻ����,��Vs���/Q�AR��N��j��i�ؘ���y�$5 c��=����aj$?���姻H��� J�"
t�S�.����}Һ��C���)��h�jjB�ӖZVR�2�3�ʳ��>/�RP������i\����Uu��j����-�6�����$S}���̓�qp����pΒ<���T:�sܸ��%L��^Ub�X²�E5��.W���Z����E5c�rK���
)����^s ڑ(��#���F�&ۇ�`�EE�/�d߫�vC�pv�R�ղͪ0�p� _� u?�w����n�~����:Pnu�룽��!{ziybN�;�/��#�ڱ[�d�c���.>�����ߌ�?!�,����y"�W{O]��q�%�8
 Q���mV�g��šQg�w6��E?�K}'܆C"��m�`�~T $� ��g�OV*E4'F[8�����^�H2�S���S�$����((��|�j��M�!�1���~h��	��툅+a�������A�٩��"��+Ɵ&��>�ϴ�̈́�4��=���~�� ,
4z�W����	��~߷�0�����~��.v7~#�si/�=��C%t�9�ӂ��?g;iXA<��d�^�Ӵ��b�ң��=��f�w�ڝE�`J��a��2��-�
r��V�E�Ԇ���n�F���pD�r�r�\���闗B�`�3��z��h��D�/(@��#`2����U����)$�;�48�"�r-��b绎Q�Tγ{�Q����CS[�đ�mA"䆀��~��˯��ǱՑ��P�:��	Ά�6��N"_ �c��E�@S�!&W�FP��@��O�kOwT��K`�rp�h��q��kh�)������|����-��}>Ni-�tpp���#��������y �.4�ۆ�D_@ɡx�E��I�chߣ���n�ٖw��4�n��J�����	���bb?�Ŏ�t�Nz�']RHPk���e��M������|f�(b�pU�sb]�n�M�R�&%��H憪+?�A�q��MF���!���G�%��j2�Ùn������"�	�H��'`2��݋����K��\�ī�¥
�}�Y�ʅ#��t��>I�SwW|��	ƞR^td�p�f4�z�o��QJ?y��OԂ(��(�BX^�U��m0��?܅R���iwշR��F�Wl�6�`EQ{!6����kW�f���Ҳ��Qw[n�M�f�Pܰ���|��د%����2=*e9�0-b�T>t��Y9��׼[yGI-%Zf�x�y��ז�.5݀
e����m��i/¤8�6U�x�J����(4fK����ȢJW�F|q䛣�C�����'0����e�+��!�S��c/DV�8���y��l��z�Ҹ��Ұi;g�a�-7�Z�f��n.�0�d
��C�����J��a����4x��-��Tpդ�8�~��H�?_���m}e�K�Y�+�������.S��0��5���e���9<u���;I�G�M��'�s���h(*�l�N���3��Ժ^w@	�3���Bp��I1sj��L�������8M	!�1v��o�i&_��U���ts*��̄>�ݓ��e�fp���h!�$3Բ�p�m��m`}��o�V5�{�U���=+R�[�Ll�J�o���ܰ��lm���\�m����fcu&0@�3����n�L��ȹ^LF�Eyou�(3��1�v� wáC_���Ďv���S�ˮ@��6��͍>)R���ܭ�j�O�/ ��
�FA0h��}������kl/�
�R>��x���\Y�|7�;):��{�m��G��I[�����޴!P����a�|�s�{�U4E�u��vL�<�+��n,����_v�R�<�3C	�)��mofȮ�VD��D x(:��T���ޕ ��BM����L�-R�$R�mL��\��-~s��g�[5������)iB��uH��g��S���p�u�w_0l�	/%1��'%W���
q*C�����i]�N�_��>�����[x����#�a��s	t��1���#7֑7]��OT�!s��Ub�i��+m�?2Ws�A���d����3����[KR"ןK�G���/ծ
j̷v_� ��kw�E�Q.\�d3Tc{�b�Z�@fc���#dt�
�?i��'	�A�
�Qv�xC�R�(�͟��2�~�3YO_��@�_f�1[��pF.�UNC9��
���hN20H��2�I���o���&����<Ykv)s^�Fy:X<M�k5)������s�&�&-6�n%Ǧo��%w(�i� ���dڽhR��'��X�.��%��bQ�}�F=�Xĺ>�T`��k���}@���Ûp�v-�'�T�Q�ݻR3�Lu.n�Sbԑ1�"�K1�Q�$�A �s�4��vJ�W��¼(d*�7�x�vǌ �x��'UMi��3dl���6`&�� �4�����.�Y��fN�%'F�Ŗ��o�5}d��;�̄y�ɩ��m�6Q�Y:����"T�f:��Pi�g2�q4wTm��k['����F;oYn̷��땚�M�M���vJ#w�Sw��������G�^W"U���Y �J�e�
����ĒӺ'����V�R�͐3vX�m3����l��v4�r���0��Lz�Ce:��������o�Ny>F�N/^������ur&��r�W3��12#��ta���P��.�����JIL�rJ5�R�q����!D, ������p'08b�������JC�������D�a(��XY���=����M�����o�PH���H��`�hi�Ϙ^;bn	ST��q<9��AC�#C��x�����Ee�u�^;���޷�mUv��?-��u����Z�1�
���,�A���N���>���&Go����Ln������wt颚���|1=���������|�����A4�V!��!�M�_�N;��>�[�n#�.p�D�8��Q|V�?Cq��fP�� <��~I	���^�-���aU,��v���<��Ajj��?Ә$SV� n�X��ϳӃۀ�kl�O%�\�f�~'<�H��sJz��q���C�h�d�1��KtD�j�Q��@��6Tz^C���������u���s'��[X~N���~����g���%���ȝkmy��̉M7&��2�ED�X��m�8
�h���9r�T�[�+��l ��b�CҠ����m�,$��:�}:��UzL'�fJ��E���7M����mԻ�Y�bZ�Hg��LVj&��:ի�»�����)�5~�����j˲�n�}��5Tގu�btb�X�+�Yz����)��m��x˅�� �R9+`n����/4�����a�8ΏXz�>�3�_��w^�m�b��}�Q�A����?�`7%]	�q�>�ٵ��q,��堯F�l^[����J#V��C*9��}�NG�e�{	;գͿQ\^�ů/�ja9���v�[��/��z���m� �1�J�x�{��D l�p:K�����1n`�ʹ�le�=���fkP�k�ͺ��� �i%4�V���+�c#&(�ı�4nCS<20�ZR3�˫�O5�ݺp��=|�I����R����y�q��u��Ei��/��$��w]��Hsh5��m(�e)�L�J��B�#l��"����� ֝��?���Yݿ�PϾ`׭�L)��H�8Y�	ɜ�j�Ȱ�џ灧0����)yed�1����#���Jqg�Xeb���,�\�_�!Q��
a�sS��T���%b�Y8��WNUha�`g�?��W\����f��.��$�X��"�'/R�gR�^��6��.���~Q����>$-�	%Xh&)3�\

Ax<{���0Q~�a�.�y��xP���A~���젡�W�8Z������$dOU����VQ�������Q�$��'~���p�D��H\$�����$ENg��͢|�/�c{m�R=�t�Ί�JZ��q��\8�6����}����4�*�:���c�kP��ؠ E�ҟ�q"����U�X�<�!ӑr�/ǌ�ۘ��K����1O��bP<�<{�,��)�V��,�V`:�Ѐ��_%2@5O�Bi�*�� �<�6����3擎+������@���=�?M�������q���	O|�r�c���߰�,�$qHN���C���)�+���K��ag�E�Cm�_�N����_�j�b�!���%D.zX�z��Y^�B��ꞍYI&}�Io�������\�|%4�R%��u�3 =�Fz_�^��b��i��ǲ�ڢ������^8�-qh� S��pX#�~��dgm�ɥ3�Ћ��>����BD$[�M��!PX�����݅��{�9r�25,����2����c�&-���p[�X>UV�l7�Ǭi�^����g��\Y����Ȗ��PF�7���V8O1�s �\"�г����B�$&sX�Զ�'88_�NF�/>}�S�B��L�R�����ۛ�H�2��?�|ז~h��L!��#�̥��0��pnEA���0�nȭ�L�^��}YX�����H������wkZ�p��QuC���/��)�����#�Y��痖��Ǳ[L�C'g��y,L��+(��rXFl�=x�z��E�Y_I�y�R��p�lթ:1,/
�DG^�x�8���l�T��õ�����)�9�/���voGf�)��m[+@�O&�8�LK������~d���Id"���9�8ʤ�ͨ��f����B,N�B�J*�瞛�s�V�vb.i�|a�^�?t�SN��A����ϛ���o��~g�C%�ܲ2=�f��
R-��4�Z����{���b�#�}
i�v.�̀�s �&�=ҩ`}��CJ�j���
b����t<?,��@�K�[���9�]X=@������Ҍ�'x�X\W�����58�#��y�16��T�}��.I�-7��"���3���r��h&���{��G{����KjO0� 0
���4�=ቩ8�翓�C��Y�Moh�S+��%<��TR���oV�V}���-1�R�>
O��O�?de�hp��I�T	ȫ���n�9z��' �߇��N0�qW9���<)�0����]9�F,o�y�X+��Z&��� N ��ʘ���X���Ŋ�Zـ��д����NG��vL7��T'MF#)��P�Q䩡w'�����qq��$� ���}�`��΄��|��П ow(�4;'�e��fzI���3Ozx:Ul'X?����j˽��>�/8���W� ���{�54S�h��尉�f�O}I�9�t����'|��0���گ?�b�\
Ⱦ����:%T��9�9�=�{�-▎	�~��͸ �2߃�^<�=�3]a�&�遃�_�W��x��uʇ[XN׹�g���i�Y��xd��6��G�{7�0���$dP�X4��E�6AZ�Pɱ�("e��[ɕyf�@�����L�ۜ����%�*_g,��٪��W�0)>@�Vo%�2�`n��l���ea�u��ࡂU@���l6��2*��E=ӻ����1zS��`�НF��iҙa��mkJ�3	e�I��f�<�ϔܧ��}�~4I�"�r���S���R��)����5��z����E��#�5})�
���N@B*1�8`�� T�Q�^`�C<��IôD~;�xQ�@h� �*f���ܞ������Gu��zfgmZ�K2+5h�:UfV}�;U11=aV/b �=�Z�8�e%�K.�/�iށ�B/:�2�H\29�Þ�AF������<���^Zv�y5nk��-E#����["�Xt���
6�RćP3�%T��d7��g��m艼�PbJ��v�xRs� �ب��c(�R<��n ^NL�K���Y�DVR�.�c�/W�~t	u\���7���N�ݤ�eNm�F�)�/�����Zk�����9��q�*�?��#)�5e菘�<�H�=Z���-؜���ǂ��B��7�Jbs3*�YCt�;�
��O�]ĵ ��QfB/)���-+<A����Z':�
>A�:��eKȸ�b�Mq&�ȡEf�`��M�J�s2+����,��+G!e�� �k�2J���#��:i�~��2�A�	%<��\�_���b�\Sf2�D��p'��O�q��+��3K���+��[����s��p��~
$�5��E����Ƃ_�-cV[mي��%0a�2���l�a~_HuB=ܢ��X�������RG	цwM^���? }����� �c�=�+�3��,�q��Z&�vU׾�-�*�Hj.����b�*0͓��ܺ͑�fy�7&hU�����H�U��a>�P6��V}9�g���D��M"��KE��+Z���&�	!�T����^�V��#ș�De�Q*/�?�1�S��0����[�/���)	�F/$�Ml�$�d�d�"�ψ����أ�4�� �M^&��h�������
�Ś�޲0m��� H���?���l+$s����L�oE�u������(ǩV�}Ҽb�2�1�+>֦vW��-k��7�ٹq�Px�E�D�f�I����7ʕc?��ׯ����@�����>��{��[u�FQj��:�J�~�������N�=�����8I߳�=J���y��ޱ��`�~}p�R"�2��Xe���/1O��*�{��X�<TeD�����ܗ��������rӂ��>[��ҷ�\�sr+�5��x��U��6k/U�A��ص�t֥��!�(W7�J1�^o�+��f��2^��r�9�:�ou-���{�B��M?��-�=��S]4��@��̚���S����?Cx��� ����*�D�П5���\��ol]��g��f�����L�Y�L�>Q�!/��Wn���$JJ��V☻��6����}W+tχ\���oSJ$LQޝ@A6B|6Ȱ����Ԝ6c�w(��J�5�#�n#� ۚ��j�uM�]�T�k���M����&_c�7!��n����0Ԃ�M����C�:p-�D�Ϯ������}|ת�?Ex ���ܚR�؟yÑ�è0 R��,��l�fٹP9���nk�
�:J4�q���7���w����$��L�����Y/�x�Q���Ql�K*K*��G7�H�m��}�ů��R�&�����Xqϻ�mjq�"��\4�W5|�|bв"��g�ꁉ��XNޑ4r8 J�Mh5�4װN.P�φ���Z���^��ɓѵZ��<I��x����,�ŵ|1x��VPдE'�kн��U�=L�ŏ���W_ ��_��a��$��/ r��K���Ѵ������˿#����m�ۼ�^�"3Ĵ|��%"T�tӠ�]9�°N�t�n_r������y�#Q����O�ԢN0S%M��\m�B��rz6@� ��i�o���@J����ؤ�� w���;�;ؾ����[n��5�>�xP�!xS��-n����i�B+�OTL����╡��;�;L.����UG:�w+�ܼ�.@�=V���@j)P�77c�l��K��&�Fy�J�Z�YenN��{���q+�kZ�����ߎQI�4i-`j��AߞY�Y5�������bT&�����x�i�����g��^ބ���e����ځ�݄�4�MF�Fș�3׿�CY%��L����߄���3]��7>�'g�1]Am3�F��`��f�8_)\ɼ�b�\�}���0������3I����O�=�\dyu^Z�%�j��E3t�L/���W�����DY�����^a{H*��P$��>��QBÿ�����m�)��\m�'�L�~�#�x�:� �U6A�dfDHԼ����J��(_z	E��{{�YH�1������rc�"Jb-Z6w �
�G ��ͼ�nl���A�mw�G�~8��`4�x.!hc��*����/2gLg��G��&�S<,v�_|��T�7������0.�4q�"�X^;� 8|��g�9K~���ޓ�c�;&�s����a_�Dޟo�����>�ϔ6x;�.��j�un��I!��'�&*��4zN��/���W�,���k"�c�H���A�D �>m�ɚ��o"�~�<OH�aR����m�ͭ�	=:-\x=�']A�k�������T� �:MS��[�s��̂��E����(v�ବN���O����`i�� ��͠@iܩ��h�#M�	���o�(���sC.a'���]iA	o�cX�a&�R\A}���N��%1a��N$�=D�<�j�l�?�p�)����>X߇��R��@z��'(B>d� ���y��F
�<�C�͌V���B�5��T�����Ӡ���;�U��o����TlÇ9i�F��Չ��c�PuL@��s�[�C����v�^//.씀����&=зra��?�1 �}�H�$���*����G��H����Ξ���}_>.�AS��G"��oh,i�ڬad�����
?�����f�s� ���xN��lٞi%l�Q��M,�|��3��+�n��޳ن;�Z�LE����"��H���T��{�>6R�ԄMI�n�1�O�C���ܕ�l�dR���h�<Q�/���q��?l���1ԟ�P.rn:�&�ciy�0_�-py8�sɍvܟY5�f�6�T^��Uȧ��wxW��)�҂�5`��9�	$�t0�N �2�F����#����L��z{y���A1�n��h5��� (����6@��&���V.F5=��gj�C��X�5���m��j�y�B��{Hh�	�`��TR�[[#m���8�`���1&�����r"0�[�NhPS�.�B��n�����f(<M��AR��Պ4�e|�m���e4�~�C1e!5R���A�KUP]V�X�鼎 '0��67�z��)DW%#B_�+E٤���2]�s��HQF	T+�G/�w+�0ԧy�.r)>[^��{koq-R_u�D7�;]���m7�սBzDp)�?�n�������m�%�� {9爁�M�mf��R��=��jA8
,�'̪(���1���{�pR���cްok�J��am�R)a�y�䗻�8i��:%'a����iέ�xr�heZd:\ڿ7�Py��|{��>z<%ʿvl�MG��!�)K�o_8[���6�D+.�8�C/5P�EP�L+�Y�ʾ����5M֚k>�����l��| �g���f�������r���C�(s�������)��Y5�S��l�hѣ��D" �4§X��UQ UG~2(+�-��N���1�˥��8�S7��X��U�9N\!�������JH��(UC$^r���s�8^+tV�P�k� ,��d�(N��XM��qdf��9G������3G��\�(8�T����c)I �h��c�`�������SӜQ�e�)��E�� =u�Me�fEW���>9���0���*�L�U��Q%{��<S���7�5ĵU��U��F��"����F����@J!�F�P�sy���Z���O�i����Tw9/��y�@?��ݴ�2*w��N^��O>�6X���t����Q	K>����1�|�B���P <�A'�v!OO ��m�(��+�CFޯ(u���c7
���[�lq������]�JAW���+��J����l�q�n7bK�>�ȡj�TFZsS�0���M�<~�1�=ɟ ��-H��JS�)7��&�A�"����P�w6�o�֟aV��
�sN����~���FF/�T>�	�I�RH�ޜL������I��d#�����t��w��߆�|�O�O4�L�c8>�ӻ�;�t]���������K(U2W��KS�_��
b�]���{6�p���g/4���rƧL��Gf��v�Z���M�{��o9&N�"����ֆM�JմL������`��JF�m� ���,�A��f�Y��;s�}F�,�E�b��z�P�A~�Xئ���.��p'��W�tM���i�e��L��
@l�Տ���+��K9@��'�b9���2gM�-&H�U��((�Mx��4H�\�;o6J�C\�N��K̈ʅ�A�PN���֪��;l$`�-�,kv�-����A��g"�(�!�²��p�id��ױ�D��ݯP�B��h��U8��͆J����;�:1�1�12w��u�-R�~�n�������)o���!;�{���,w�yy<�V@Yq$���ļ^`�Om�7�<�|5p�?���s�m{�OV�h�J.��Kd!<�MDHH�Y4��5����`�:gB��&�҃]#�D����]��ѵ�3�_(����L���rRT|���X��Wen{%'�U��;6��5o��O �.�Ҝ���y>�KvE����~&r��q����Lי t&v�P^���j	W�6}g��t�u��؈�O��/�����0��@�J"
{�Bs����{�nv��i��Μ�4ZPC�7V_�]�H� >�؁�V�lq�gX�0��$|��=�
��p;98<���R�M�q(�F�ѕj?������?�Am���a�@J]���ŖX�Ũ����@��d��q��c�F+�q3��j�Oqᢡ�[�6x��w��]��c&��zǿ�� ?m�;t
]Y���@�d�H40T��?�EX�P�yA�@f�ab�h_���t���0o�7Lr�q�V� B���)���j����+�m��=�~<��� ��@�mx��ĵ��F��#V�G����܈��X��SGn.�"ɉ��(�@�S N�V"TnT���1�ٖ���� �GK�h�nS��!? K�jm��9���2���q�Ơ����vY,�ӡ.KR��k����V} Ij	���;c9��^�B�Y3�� C'�fF]]����S���(��ӂMp��f��#���I�<�y�+Ak�M����&*�Z�T�����7�E�;(�s�jX�<���@`"(x���m��v�)2 ��%'�aQB�Ub(i9�@_�ూ��(���obЉo�k��uB�l�ŭ(���F�q �屏fe�w��3 ��c��_hm[� <,W�?a��ACQ,̥ '��M>4^���j���XW3���}�ZL'�{�՛
G����AH�jʆ�����"!
1�/���2�:��tS���y��:�/��nP�-;NЏ@Гl��9$5o	�F���)fQ��C/z	 ��t�3b:3�Eƞ�:8�#���#��ћ�� �(�b��<�|�<��!����EY��	`�y�	E��E�{��
��<�x%��tӑMx6EZb��4g�c?�qv�!�s�%A�y�<��[ݣg��V�q ���M|T
����Y�L�K�F�����H�D�)�:o����R�3ي@'0�L�d'�{�ȯ�]�2���\��OڬK�sA�ѧʁ��rdIԖ��P�W��HJ��������?��W��L�jE��G&W�k�Q�ƭ�ޞV��Z�E]N�>	7xb�S�^h�O���h�4Ak��m:��7���TH����=Uw�/'�F T���&a��`���b�|�w`r�(�:+c�!2��ka@�n�BG�B��0u�.��NJݓ�l�Ш�T�uiȫץ!���0�1������#��6�[��$+���dZ�FF_��{�g�HT,g��Ζy�'�4�o�,����Hln�I�-�V^r4V��������{,�(N�춿wHt���Z"X��¸��|/y�'�E|��3c�?���z#�JÂ�1ߤ��Vj���uH�J�j�2�:F�T��zO��9(�m7��6��p�������i.��1��\�2B=�2E�9�([��z��>,�a���|���d4�2X�?���g�hFS�����IZ�g�Q�S@^Pe� �C���"O4��yæY�@��.v��青��CL�Ek�]��ۮ���$c��sE}�[.d�g�zo�"i��g���Պ��WIp�L�����gX��a����v�d�7y�'�=�r)�!�QG���o��<���i��V�1�kN� 2ŘH=�i3h��:����138mQH�X�w�W���ʭ,��9�@���i���f��3��{'��	6T`�#}%�E�0�����5hʣȃ����W(�y�;ԍ.�PP�_��$���J�����h4lcw�F+��� l�G�O�����g�S,�>-Ȓ��1R�兀�R<���-�fȺ�����W�/n�f����4��f�rqNR3p�Ĉ_�SFە\�l��;��J��5��ߢ��P�X�eޣ06�`^#� ��c"�EO�lɤIwG�#�4�1�$,{3#g���M���N���<udCש�{�QW�T�ɺ����G-�W�P;��e�ࡦ����� D����B����a�Y����F�T��V�׀����P��Q�l�XM�`��µ(���&㫬�q���88o��:�kv�6 �;~��m��b4l|�ZN"�-uQ�T�3o�����v���";"� nB�M<h��jiӖ��9��2��Cϗ��	1��̷	%��b�^Z Y�N)����+|�ׂ  aQ�p���P�g ���_n���f�994��=/��_o���kK��1(���I����O*���V$�<b�8��aisq�'�DY�wԤ�'m�؍��Eҙcp�`�42��G����m�{�E�x��<�tlې��
�z��|n�y{dkD�c���~Z�T�>�2h��XK���V�y%X�٤�vu�>�p��L�Vp�b'�̐�<!�L^�� C���aÌ<�J�h�+4}���I2�*�YX\� �NP4��E!$�G;R�g�Eq�S���+��~s�B/�(�-߲S�r@!���,�z&gn;��gI�ߦ�.m��w<�������+����/^
|�� #/�F�[�}RC�[_Qt�V��'��D��ps
 �����xͷ�����<�(W�}
:캤�ZH)��Kt��3�]���_,�Q:��z�sh`Ӕ�#��~6��M�o�&�v0�Sh�D�A�$ �U��D[ѻ��b������lf��h�k�W,[��.Yض=��z��-���u���%��mԬ�0�ǆ&dw.4zQ��z��ZUBuwD����9m���J!�&�⒗�f������� (�@�,�[�nd�q�`��k4d:Ū�_�C�	u�:��4O�[~��v��e�ӑ�`>},ƆL�v<-7�+���������^�C������\f#m�VEnh�E59%��r��*���"⎲��nCn�D<�6#,��
f�¿0N�Gn�鼞�����դ(�g(�jzet��,UC~G`�#���^;"]Z���
�W{A�dG+Ĩ��Th<������?����r�#�4b(&��Mo�\6�8}��K�������B|���'<+r�1fk�4U=귟�8����Q�x �>]�4M1�e����Ch�Zۗ7AȆ�;Q�H�S��0�_�+����G�x`�~>%/_J�u�eM���o΢i��v��U�(�c�Qd�8
6��u	�6�辳[Rl
�.��`�Y'k�;����N_�ݾ�y���&��x�xn��x��
)���Rfw�d6o'��v%K�H��s���ͩUP�|ƌ~AͣrP�i/��"��KM� �J��l��f莿?�f�oCS⤖v{w�����b��1��ӓ 茢�g��4�-����I'��^���p�kD���~���yAB㼀�3U�>�Y���d�WE ��-����ͣ�>��VOƫDESj�����8qO��	��v�ؤ�JzF��E����K�Eղ[�v��u���-���{W�tnm9�l����B�b�j��t"1C���̴nm��
�dȂae7�!���%�xH�V�
�X�l�A�7��V8��c�2G�y/��;t���t��/�m��a��Qt�Q��{�d���s�M�&��<QxpW5�Ð�뙝8�B�Pc1Rͷ+�_�~��v��ƭ@r鬈cs�͛d�u���G���l��(��k���/����/n�5V/d'l�5��S�� qjDΣ�x��G��oL��B��E�^6�sp��rT���,h��T>+��l�2���Ǔb�m��{d�k�p��������1Q������'�3vAg�%Xz��DD��#�\�8�WjT[y\?�����#�0C�u�oxz���Njqׂ"�C��zVEfDt�sqBGzҒ�(�v2�vO$Ʋ̚b��"a��6*��?��e��;�p�Rd���HtA�������Ұ|���Q���Lb
���w(_\�"+�-�	�0�X"�̐�a���Q��������F�3��ӹj]����4�����$ALC^����� F���Q ?����}�N��^SU�a���{]fҶ��@JL�k�Z�+*]����ZDx����s]C�~q�TR�O��gS &<�1��Y����;�v����a��m���0O�Zu	J��%���}͙�Ь{W9�;�I��"�{��ҥ���E=L0�>�4�3�@g��!�A���\ m��.0=��-�ʳ���%+E
0ԃ(�>M�1�_��Ȭ^����xz�cp�[����|��O�i��-蘊 ����8l��z���˷����j�c��>����r4tI,S�/)������6�%���}d��9�ؒC����RĤ��~�%�ڑ{M���Ȏ ��Yʌ�� ��H4�o;�a�/௩D��IΘ�ZAA�J��BL��w5c�@!6_K:��+�;��H�7���2�g�����ȸ�"?����[�I�)6�{��v�˪l5����J��]�J3i)c�5��9әZ9��}>��0����Z��⤺u�T��B�S7�a��H�Ae�4��EƵd� �|����y���B�|�Xc����^�:G<��i�JP1-�Q��/��Qx䅜�h�r���7C�"r(��%q?Ÿ��x�k�Q�����혼�5�~��,ޘހWhD�(t圥�RAs�TKH� 9����_H����[^�$������$�����0��^�<}5>*ݜ��w0E"����w���2���0�@*���	�M�0��ӥ�hzft5��~���"(ħ_�W��{<2X5Z|'�@�!��/cvr��N�oe���vk����,�?�^�]���}�+B6���1��u����$�	�\	��
�Qڢ��0��\�`��[��6-��8��9��p�	��Flo(1u�.D�NW�=�"Wv��fK5��$�~�.kA�T��G����ǭ��fjN�%���B��J�f�ܷ2Lx���$/�%�)��+*n������t�
e���dt�(���iF�M�!2 
�U������^���\�em��ӽbuB��,�Φȇ
�Tp���Qu���M���Xvȵ�G[�TC63���p,���aF���{M&���K�^�J��]���Ǣ+hr�ܜ߽O�ɒf�?­S��V"�{��P�����2V�H��.�,�JZ��资����i��ބ|̉\>�
�S�&=$����}BJ�?�
"�M��)���L��qt�W!��YU�#��t�᷸@�B�oZ�' �ަ���E+��S����.�����eIl8/��!��.�7&Oo�_w��d@���Ȕo�j�/T;�m��YӦ�tE��7��4^�Y�ћ|�JJ9�[���Sh�=ߊ��y��:_	�o~���Y1����SM�K��I\P��V��K�#H���Q����(8H���΃�br�g��S9Z����:��Q*@&�%�A�(��7�7�s����<'����<c畉t�Z5ݐO�/��~�cb'"u-�SQ�w��ǥ��u��|��w1lU6�@܇���3�ŧ�������܋a��e�_h7=u��sKtC�F��g�](�qNv�jm��G��]<{�y����0��Q��4����{0;@bj��`�T\�2[�
%��N���?6a9��-T�/Ԭ؇	��'��KB�˛N��\{���-�x�>�QT�So���'ZO��jS*��sYn���lh��� � k�'�<�$ȵ�ļ�-p��{17K���)��^d~00�:�ZYzq�1�0�<�Df���\B~j_�z���"j,�D���|���$�J��z�v�n�!�(B�4�<��VG�$��ɎY; �%�'Q���Ԡ�)x�f�����nTd��z��'d��d�ϧ����&���Gj�R?C�f`q�cVt&~���t%����U�x�k���m�.�Q%۠x���wƕ�f���|�A�#��:��m��;^}e-�;���lAcz� ����&�P��A A�vᙙ��U>�� ��+�}�`Vp�{)����㶿a���s����$�Afa� N[3Ұ����0�Q��߃S߂�#>U�i	>���z�O�ebv?�(3����)xw���ߚcV/XR��"Op��^)���)��T�!~�)W��NJ���� "���t�r�A0�-�
��Y�}�9.��o���$�"��H4�{���?�Qo��<=��o��u����FcY��+��w1/�t������ɩ`+�Ӹ<P��
�Y�5���nT{�	��r;��|{���V � ���o�	�\��en���n=�7���r�껌$Z���,Q�eQ�A�@��	$�ܤ��=E4��N�G4��I�l�BN&�,�5�m�Q��`dI�z[s+A��e#5���[���İ[�;@�V�`k��Ób^�:��E���|(;�0�>�CDv�_IҤ��'ˆ�R����# �6lX��I�V�k���ੁ��[*/��������EǨvh����;���!1���b������X]�6���;��P��ԋ�f�Z��Mi)���?�*�/��n�k%���ݵ�����w�%|�e�2�}ͰX�u���K��b���ƝJA��_��_���]��6izٽ���ݐцQ�uRI)B�i��n2�������!
��x����-�"�&��e
��`�2#]E�Kh�s�G�srE�6��&������j�n	�u	n<. �5�Ǘ�)0W�ӏT;����/x���4�J��We;{hS�|����9����(�� &؅!���aJ�z뽃��)�70����	LӆL��_����$���"P��#����
+Uh��L
z�h���m��W�cmd�{9QF��艚��yיtL��,�&>a��#N�6;AF`1C����m���
߯?�~M�	���p�4�I_���g����b +"����wm-���l��2 �6ܯ|�>��y\��Z�NU|��a��6���);��K���O�Mۨ�$�8o��jA���(`[�NF��T*�9璟�uR���a"$L������5�X?�+���%��}GB��j n9be�������B���g�^߭:,��+�YŠ�Dbu�!�=��,�����v�^�ʎ���������c��6YkZ_
�O��(*T�f����+^F �s\)�0r�F�o��\F�����l�	\m1$5Y�������VX����G�V�+3���� 0Ǌ�h������Pq;��u��z�	�F ]J�������X;�!S�'���o!��f�,C&h���[/�G��d\�+��,�C��wU��ݜ��c
��-|ע�ζ��d!_�%�wR�.P��#�q�z�Њ�p	sA7�G�^?~.����r*�����[X�n#]��tʁ�}���oVA�~�iЃӪ^���z��)��Z���
�;-Q?���!j��l=��c�u8�w�j��`�ؙ*�ʲR��o��>p��N߳y�>#���.^�B�
�G;��8c�:�eǡ���2��$+]v�Qf��?n_l Ќ���hQ�dM$ KbY\M*9ܾ]�놇PXN��_�[�EF�L����<a�k$,�Ҝ�Z�OJ�\I�By9v-ىO�>�P����xnޙ�gyu�]�[u�4�xt������z������?@=�`^��I-�������3u@��]|6}��~�C��_!1BE�(efН�F�A3���y���UBޓ-���M�9P�A[�xo�hO�m���8؜c�wH�Y���An�0C[a��Mɉ. OE`��TI��?��:KV��8Kё
3m�
;�Bi�l��}ȷj^��C�T���_�lQ�T���WN�&���_�SJlg�I�\��L*�Syxs�ĮeW��=�ʟUaX4N�V��긚�{Խ�gSo�%��C��`Ŭ�N-*��v�-�a���-�������/oy8#����Q �Aa|�J��y���zәW0�pxt��+�y�C��[G��M=.O�$�X1��1��$�
� S�޳�tpjY��^ё�QH�mܪ)���2�Q�E����4���J�]���A���~�|=�����
��#+޷���5=+�LX�6�'!�1�D���ܓea����S����ُN�.y�� �\�o������hn ��>u%��CE[�f&���#K�c{��5���4�X:�b�R�f���>A���ߒ���>jU�ȋ���x	b�Qw�[^Ş��{@n��V�� �w�a����-y
�|�����q�~-�8��N��)� �K�^�g��z�Afy8������1G����"�<l�~�Ǵ�����'����y���(	[J��Zl�9H����w-v�J�5��D�pZ��8��lj�k��Z\��Q�����$\��a8ǐ��H��np�	ĽMR�,���$�-�ڶ�J��!��An�\���J���;�I�� T�e� j��̔k P�+��,	�4�P�|�j����-$��ҡ�:�eR��P�\�H<���X)0�@	�1�4<���U	�C��"�8G������w�����s���(LC�v���ZO��zS��?���ǧݿ�����%O����[�)Iy�0D�x{�~�B���6�^X*|�)��C����vn��������|'�M�#��;�gj.1a��߬��=i��6���4U�w/�ȗ��`����ؼy^�Q'������	�)�cIR~��%�sҁe�":�Ñ�ֵ�K�G��;.��u���sT�=�J�6M*�A�����d�G�h��
/>��x��U�
z�~b	@T Y噢 0E�I0j���.���[mC؀�D��(�wk*oU�Z��[�_�bJ��Y΄̭ �ol��I���w��nu?6M�"�.=�ꬆ3���(�+������&�;������u�^�t�Ʌ�IE�t{�U�6l5�k�=벝���>�Z.�hq3#Bφ�`a�S"�󑓥��$O�Xi��jP��N�6r�8j�:R&���at'��a���	� �c��j����z��n�kSxS�{�DY��H�X����DFXu������W��д
%~�&N�)�r�ڽ45:?�qq�A����=)�9m�pLr(��Yh�!DX�p���M�d��a��m't��l5�V�Y'wW�����^$A��c��ok�����̮��$|�ZhGd1T�F��~�M�He_B�bvw;�/F.ϗ���T��V�j�#>��z7 !�)~ݖ�G%���p�8i�3�	m=�H��$�v����=���8��3"���+�w�� �H� ����r�S�z�E]ɣ��F���h�20),��v����Ll���>�L��������b��J��'$�<ڰs[�`Q�|�ӆ֯皷H�t���UT�L��b+�{u{v�`����z0��%��>r�Tx��rD�{�&�r�0�h}%N.�M%*�/Y׼/���i�r��{B��⾽��;������VB�j��a�2G �GG��E9e1It���#��/X\^����U�%��'�=c��͠OK3S3p���:9� �a_��[�g� �
wy��EL��"��O1� a����
��mU�u�ѽ��d�l�Q�aB�x���*32K�TC�@o��xn��a�AW�g��!_���*`�
P�0�iy�_$�jWW;����:pNբ���2��ޙ�Ho��wV%�O�C�0�?:���'i��Q�>I}���ƾ��g�>KC��(���M�2R���:;[�f�7]<���8ԟ���L,�Nx�m�;����:nt��ӭE.R��/נ'��Rc�%I�$2���{��<i���,��ͥ��EI�0�8�8G;N9�TNL��ݛ����V�e[�jׇO;qy$�@b�#�I����9��}��S�}�㮇?kA%s���n�`��
�+��6}�D���k�K��բ�$i���ׇs�b��sd�6'1{H������6�j_T�;�#ڂX�K��<^M�f���_U��#�ٰ=OM6���5�Y�R3vG/����߲s�/f���'��w����Ǹ/߬`'�����a��RM���
�f�t�7z~mWB��/.ks��)������?DJ�2�z"�ES��Q������ٵ�Y|�omlg4!j�`W� ��tq�kM�k��_b�q�	��52��1���]̨�H>@�ĝI�E�h��?*7h�{&{�>y`X���o1In `5���g+v?��@�s��\��j�,�S����l�����ɼ�<^P�0+*�4y���(��E��r̭�'Z�� 2y>�����Q6��D��`��p��{�]�g��.�*[v��'�;3��>v)��	3w��
DI�g`q��8���L��^���������H�������ֹ5_ղ^X%��O�>�+��nu!�ZbV�.qX����}m����:Oa��,c������|@fC
�c'ȿ�pϕ���lF��juG��9���Ć2�;_���߸��F��*���P 8|8�O�Z]�m�$x�(qnY�y��>�~���1׊�I�K0��7$*���2iA1+�+��61������9	&9W���'�����=�>�h�D5h�8ܻ=�1J�o�yG�%	c�{�m�0��~��g����S)�|A���<v0���qF7d��W�(5`�m0ǧ[Hw~~*�m�#��s��B�En�Ѯ�]��﷑q7.���?]4�[��Ee��#�ƌG��!�	Y�/���[rW��U�қ�vP,>�� :�Z!��L>�R�X.i�p�\������k�0�-�
�Rvml�I��C����f{�ۨ?�??+r�sHP.��(]|�ɦ�\�S�(V�e������w\p�����0��f�� ���܌�M?�RP�:�g�Έ��"Q�U�1̘�H(m��؇+��:^xr�\��`���*cM��qA���F>���Ex���ZפU�Ng��6lAcMy��ߜ�[��������}���q�#�j7��Ԩk.XRW�j���c��ۄ٩�|�J�ؠݷ��J�G��4ȮoZ�fvh�?��s
KpNK3Y�n�{���U��D�{�~�u|h�h�ⶏ��=�xy���X'<v)�*�G�x]D�z�{�_�@�-[�����X�3�o&A��$�C���*�v�/D�&�5�Y9���n�o��x9���-��R��$}�Mٲ7E)�#��NFY��rR(X+����$��u'M��Eln����/���[�PTv"���%�.��0:6�� tf}?+L�?:H?����J>�&O9;�
���i���I�ܭ��lԞ�-�"�Q��ɲ�2��b�̓��?u����r���m�T\�����G�;.�r�$����ݒ� �L�SZ2��c���`������ʖ!|)H���H��e��ʼY�wV��8'����h5���p$u��}�����P�t�ϬW���<bҎ��6��p#=),��S���n��l�ś�d��9���x��Q��.�e���{�@��JHh�rOd%uD�e�4kXĞ4ߧ
��J�K+P��<ma��`"�.��d��Q��a=�c2H�'A`���5�vԶ0[V��t�Tb�?�����B?�G"���PNaJ��H�q^�b^N{,R�R���Y��R���B����4��z�q�y{� ���o�-�����
תS�w�5���>�7����B.2娡#���W�OD�CZl����艖i6��BP��]��͑N�'�{;l��}"�>�ՇM�Z���~0�P>&_��WC5'�q�|_��!��.�I�Xwj;�a��9���I�1�h�r��p?Z�u�������>�q�=�`�EG1��r�,�)�PkC�N(���ۚ$�|A�1�TU�z��%C31��Ţ���"Ɉ�q�:�HJd/�p��Fm��q�*N�چ�1��m̺֖M�1-�wO��VU}�ħ��y�2e߼%�w�^�5xMb���1~!�j��SH"i�m��r2'�����wȶ�掼�=�}<������s�Q���q��}t;Q�HVy�b�-F�o�x��TհiJXbh4� I��N�/�����v��T��|��%���K��/�ϠB'������>��r�,��^{A8�U���Jl7�4Dp,Ai7S��'(�@�O,Q٣L��o���lP��Z���[x����{	���+��/�iQ'�[����BUi�Mbib�?�un(s��:R��0~�H��̐���[�R���S���,#��֖/�l�A�w�v�%C�ȇ��v-����s��s��R����9��T�xA�_Z�q��@�G	F�W��D�(/�rj�	�[��"�]j�|��@�Bai���k<!`?�L��+�.�@[:{zʧ�<q)j�SY>��/�_��8�sw�!�e.>�UX��}Řt�b@�e�U��,�8ê��*3_�ꏪ�~�V �H7�e>vo�#��<=�������%�P�aMS�s�e) �=���a�5�o��Y��W;Q�I�7P���O���fFpRd��g���͎B��y��-
(�A
�'���c\f��T�J$~����5����u��
y�޳V� O��/�;+l�k��gu��d�ێ�$�ڑ(I:��4%�-�)�EI��߫�
����٪��h]M���r�l��9�Ss-ɗy��-><�GҜ�yofyLXq�lZ�{�o`4�㌴,�Ŋ���hN�1/;"~�)���G6A�J�L?�<|q�Siv�Co�0�δ%'6�]�?��R{)��k�{���
�(G �����2=ւ<˞����o͘�w� �]��:��;|K�ϙ��%�@��h�a��)RQ�&�?��Uf�1���2-Eq���eؖp���.J���9xeA�i����}����3b�(`y�¬,��d�2LGi2V��%�XZ���b��S�Z�X�/�~��h����'�����V+R���Ĝ�*V����O�"��![��(�1�d'���n�[��8��ˢZ�f��xX��).T���@j	��mic*Ѣ��T�rw^?	��7�	��,{�C��2F��Yx��q{BXeM��*N���wv?��x�@q�qֻ���o7u���fP�v맷��G,VK�H-"��;ٚaJ��[(�t���_��MG	=&�2@:�����
��)?Lh�Q%Z�E� 3�+wn(�����v4F���a���!�S}���f�<��Dh�2H�#���a�X��oU�ȍ��J��AR���n�-�[}�f `)ņt�Y&�"�g1�����t]��%z�@���oڡ5l������C��q� �n����oȴ�c��Vc�Ya}V����J�a-݁��|�ۭ��͒_{��|?�roԼ7ؘRb#�T�Av8���fgsc�~�}���\�y�a�ˠ�RQױ�����:>��I��6tѡhx$C{�Npx��*iݚ���2�������� � B�pV��Q�a�����7�"�*h���Ww�r2��ᕂ!�i�,�vz�F��B-��2i�6s�� ���%	���!ѕ%��}���m�r4/��ż� ��t��甍�p���l���v��z���bd[��=��pD��ySX��%��8OД�q���w�T��3�I��l�:a�_Gd�=>����d} 8Q:0�D"���tͻ%x�;��"e /`�^�OH,Z�y��[_��A%�,��+e���65	C�P#�߄`��R��w�vӇ�pOE�AĔAoc���p�I�Q�"����	ݨ�k��+�y���2󧬃�#(�iF�?�Z��a �i+�o��Bt�Sތ��;l��Ql����w�I��Y�pP��I�x${��PR��� 9ՃD��PX�]�y5�}�����<�N��҆�L�|� ��W5�3�E�rt�)ϲ9����ٖ1#��O
�:�2��q4g�h�������\���1��W�I߭�/���.`f�$Ȩ��xE�ԌpKHA_�{Pd�:{���'�n�X��Gs���	�s�7���ͤR�*��(Xiq�V.��?�Z&�����D;�m��bRh��#�PE��ܶ�.�ۄPg@��ی��#9���w��R�T/š�F� p�p����p�0��peF��91�I_�]���ԉ%^���~�,�C�,dT)鷵���G�o��6�9>�i��8��? ���m�c�s$�bfs�<R۪���  �£�=|����:�aLg���Ƚ��6i�~}��؉[���<���4�x��fw�>1y�F���<c�) �Cp��/����<���.P�S0�^�ڇT�g��z�3'��
��R�i��OK�F&z�e]a��`4��g��0�㰳�^�?��T}-�J����ޟ]���*�����a ���&�F���Q��>.�P��C_�%��+Y�! E
y$f���Q�ΡF�:ɨ�.�&���b�-+ �Ev�E�o��VP�Њ�YN��.��Ӆ����M�KQE� o�����	���T���AA��4&�����_���i���5�MCg�6h�]A�� �ZI�6�Qʩ��Q���@H�?4�@�/؉4`f���U��K�,L��1���Oǩ�٣dso��r�3���3����s 	���{ 4P={{Cu��U`|����\�fM��aSN���dC���S7�� �v�w��h&	ퟤ���?%��ƭ�&�oKV��g�f.7��X_�f���.vFpq?ڹ����ſ��Wa�s�B��v9�q&�"Pb`s�`b����Z��	ם�+8%|�>���U3�l���.�ӯX�a&o����+n�ר	�>�WkN"v�5�e+�$4�l��-6���I"?��5���`X*K��[�&�1[hn9 W�o��5Iof�;�ı�6�s|5{��]&?a*VT4e		��봓3V,3z���7~!�d�F��DS�q"8�)-T���+�P���M�E����֑\�Zn��+P��,�?�ßc���L�e�l��F�ق�:s�.�N[��	1D��VX�0q��*��6�a�۪l��.���"�ΌQ#v�|;yIU�y�G�y�둯a	j������_��Y2�Ǎ�*C'L��qw�@ ��|$S5�?��#@f����S�u�fvNH���k�bDAT�L�����D�c#<<V5#��}�<-ҵP*�V� 2��'����E�8 �gP���H��a� B8~��'����N��3��;��>�v۸ޱz����$^#�)��D�i� ��Q�ن:8�~�혏��^p	�ބy����܀2�1B���|���zn�?�1k�A��:XʷRpʗ`�T��բ����Z1�nޘ��n �3��O2��ؽp]!�I��V+�e2q������k%sUL�!܎���j �\+_�B�ɯ9�>$|������j���"����p���i���Ӡ<
p�DԢ�<`�v�_u�������9}�R_���5|/����f.8Q��ye��ٞ�Ċ�rL˞Ҋ?�[�#/��;R�l���|r����R]���X���B�d���ͤ�4|�;�%�h�Hdr�� �7�+s��i^, �ʽ��Z����Me,OO��!�E�Q}�).���r{��B^2y�jMa��=	�8,��Q�/bW�����E�H�K	��	���yN��/L�g?��N���x����z�#���|L�^`O�[ )��Q=wE؆������E�5�ޝ���(x��@�t-�;����8A�a�Ԝ�_Լ�({���h\	ň�%�~'�ZB�G�AZ,r/K��r�O�Z��Z����I��]ʛ�b�	K�G6��1������L���#�[����ϐv�C�u�d���7f1��G�B����XW����''ålSi����25�g5�����71J�C��P�ʲ^(�죺�ð6ZzF����6D%{A1 y����i&�f�F�u��>5x2Y.�GxeK�>�{�*m��x\�@r��F�h��̧XW�GZ�T�m�p5�ޜ$5� ~��FM���q�ا)Őj����_��V��-EWM�hm7�ˀ<v���Z/�5���)Y�ϼ�e1�[�x�}{�U�ƛi0Nr��Ȋ��sȪ�(�N+3� ǝB?*ԋ�z���w��U`��5���y���l��V��'
�" �}[:fى+pY%�HeQ?��=ux:����R�0��r�V1�'�c�*��S����얛��BT"+o�����e�-���Vrw�H�P���DhnÈ�M�j��d��:,��}(<�E�c�y� ���)����ێ݂�g���1R�Ht>'��s�|C���ogs��m�a�k��^�|�A�������`�����O��b��R�
{0�����/N�+���RYYT�	6�~[����ߤ��(LkK�3 U���şh0��@���&UY_�Nz� ��	D�;��\���ӯ��ח�l#.���M^�T,thJ�N8�px4]�R���÷8e���	�2jw�?�O����k%��b�1�L�.`%Q1c1��x��
�9T�!k�d�Q$_�^K�2���xPu�bJ��(�����FQi��ꈉ���o����ǈ8z*���3�)N�-ԃv�DIs���~h�F�/0Q���M�i	EͰ��L��j�]��n�噜; �Y�-��a��f�����2��Ӌ��h&���h�� e�p߭I�r���g���u�ly���|"M)U����,1\��{�#�;�o���=��������jau%�x�I1�1���i��c}���'���ˢ�L�p�������B���!i�fͤ�c�M0رȆ$��a@4�
ot�yjQ_؃[Ԃ���ճIT_>D���=��7�8ڿ]�ʶ3��>�s��=!�J3e�U�\@V�����[׸��J�<���l`5������P-"��%�[�it�)(Ae=��\G@dh~qF�?z�'��Ѹ�cJ�'���^��Ҷ�`�~�k^����w��j�ꍪQ�~�X�a8��DAѴ��W�%'F���	D #Ԅ�:I/�&熩m�ˌ�����L�0�7�(�	����|jnf���73��Y��rR)���8��&�}M����p�'+�Vi����2r��m؎�,�6ey��G��R�h��	�\�rȾ	�x�һ�
C Ͽ���I'�e�o����κ\��#r��pN89�#�ӏJV�� V
�Q��]r蚹���Wi� ��>�k���lz|�rPP�IVc��cm�H)����m���7��*���8���e�'��y�B�rAC3��u&������G���u�( n_/���RʹU��,޴<��H��J!�R�} ��]�;�i�[��9!�X����rbf�~�R˳Wa�O�
��&���j#�d>,�(P��]�
���*²�����[���"[ �?��e�i(���fn8Zz�`�6(|t�,���������Ot>Zk�8Hjv���l��@��'M��LYʡ?�ÉZ���JnO3&�׾�-�a�d�k,�F����+b����O)$%���b/���<�f��5�P�)�9��d�k���gO1N������)foM+�/3JE3�XU�$:�i���lOۭa �i.�����<z��P8�9��}o;SB�À�hu$-�p�����7{�+��M�F+x�k���2>�A�C-;Y��FE�[��z�BL�|[,㖶Z<�a�F�Sk	�W��F{��F�2�|���H�6��l��� ����}ՙ�D��i�h��l|���c���_3t�e/��8�'���g��9�D�Db�/��V���σ��4 �:����&�[v<�[�x��$��EH�j�JF�������]��h�N���ڰ������+ȁ�\*ׯu��%�A
�)d�Ug�s1T���eh�/�>�g�+_���t�ceo�:�{�$?:��4_��s�}v�EY�P�Y��J76JKHޡ���BCa��}R����@�#K�lG��ѝq�IT�<��)�����C}Q��|�� OZ���km��x��t�7٧e�>�KX2x�^��n��|u:��7y��+-�G�D��CA�c`
�"QüN2��
!�C��'�?�i77�Oz�J:�M	�fFf^VOHo8�/�%��?���&B�E�|�b FDm{/%5�h%�Z=&�{��(/m)��8���8"&9V���$PpYPu�aI8 �+�,*2�iu��|�e��zصy�F
_.Y��~�< ���n��9U+�v�G�Q������8cO�~ԓa��B�ϤfP/Y�!('E�>2qb`/Zά\��=�N=GK�̟>�lHS��� �*O4	A��2��.���
�>SfUr:�b��q�K��H�YJ�̎�!�v؉0u�s],x|�����Է{'���k����J����ș�.(�G����x������6 ϝ%ar���k.-�����i�^u	��i�y'-0�u2������e%Q��<�A������71ӎ0�b�������jQ��ve݂�w5��ԕ��[ۍ
Bzi�^�Gj�j��In.��=�Q5C�}�P��*���q&���\yx�7ܯ�R��Z�¿��M��2�Q�m��BLޤw��J5���~DZ�9��5��7��*!9S%�F�Xz�b� ��7aX���ԅE�ټ�0N��h��QPE5�8��|e��h�f!���a^�e8ݗ��>�.P�����Ōpֵ�cw`#3_5��j�Sb-��� ��TǈC��y��,v�F�Q���m(yC\���F��h�&\3@� ��VEz���͛eh���7��!mŝQD��}	ڿYz�
=�h<M~�CI�a/���,3�W�ݺԶ!��ھ��V,(���cEaM9�N7,� �<��`x�F�0\4uLw��v�����/cF4`�ց�����W�E�.�WLF�� lo����4�8DW�6z1L��\{.7l�@,��
a ,�wb�Q�$M��X���7��朋�F���� ��Fw�Q��Cu��kk�DQ,�	��^�^4�X��Z S{ P�ȣ8U��5�-�R�N�^E`�`�F4O�鸂��Q-��nS�Y���y��|�������򅯡O�X�UrS��9]��!4���< %�Ԡ���[��)���4� ȵ�F����R�^	����}�ޡ�[z����l	��CC�J�ox��,��������^�
����hjԘ:�Қ��`��\���?���X�wWX��f`�Q*"o�Ozk���\ʺ&C��1��{�#o�A=@�T�xtd�,���)`���qC�ubo����E#ٴA��k��u}6�*k3��b#�Z�(� �s_V'^���V����G:�ƞ<��5Hu�ϥz�[������
�����y�,��,�t�C8_b<x��%�mVԭv��t�\W�j]�M��'��9�~��ë3����7�%��ra�}�˼�z^(l�ԃ�f�?�z��[)�jr9��v�!���$t�,�-�֊Y��!��4��@gue��H�%j�B����<
/��Z%"�'8\M��^���n�-Ƶr�B��,�ux�����)/z
����|QKl͂Z#^C�X������G!���V83���&a�/3z���@mz�%��i7C��.38SkL�뮞�,����zҢr5���u(��ks%0vJ%��O�����E�*��d��lmp�C^�W�j�)��%wJsO�
}����!'9g�|�w^�0��+��ꀜ��犥e�*'��@�o�!�2i��+��]m3�'��>>����e��d��"��u%W6=i�';;惡U�� �s/7��̿��	�WL�iRm�l�?�����?c����Q]G�������I6���3�|�G���a5,�����o߶�~�ŀv��I�P<����0G�
���NhX�L0N�:�y�d�d�
Z��������G�CB������V���n��"�'�cҒ���R6\�u��m|���8�_d��z���%~�0K��3 s���~�w�k #�f;A��w,D�#m�X��5��:<��`��}D�z�¦�GF��b����3g�����Ϥ&�Ѱ:�NgO�q��A���hs��������s������!�� �_�����B�~��d˺�cL�i���y����>��JԪg� �B�V�T5
��9AJ����cT�I�����7R�&�d�?g���V�E������7�U+_Ȱ����29���n/�Z�J{�>��@尓�t�DUrX����
��ۍ���#�.J=;��AlW��h�'�-2[�gU(�A]d��4ܨ����j��v��	��Հ�9b�d)������z9l��(��)(k��NW�����[r~�WT��-r�z*�iJ$��I�˽��w[w��g�т�3MT~y�2�98,�<*&N
��0<�lr�a�	�M��t!_������{d!D`EN�)t�����WA�'���2?T9?{�5'tXJ�5�}1[|���f8�
MGP�Y���$hq��S�J�\�w�D�>�J�{�J��>�l#���Y_���e�4 �h�|����7�)^��k�� Y�{�]��sa�O�M�n#<C�Zd`�wv�+��^��$�џ�	y��6r�.�A��kci�2�^ 7z"Ҿ���1U�ԢTʢ�������1v~��ms�~]����-��RvV�7&���?�\5�E��jF�i�Lual�|�07�]ypR��R|�:�Ϻӝ�� Jҡ��U��v��:(4g_y�l�Η�,� 63v뽩Q+Q��v�ے��ё��|WOd�V9��X��Q������B�4IUG���ɸUN��Ub�ހ�0�t����E��TtS�Զt�s�l>ņ&�d�n�o��P�.�ڌ����¶�Q������i�*P�;���C�A��a��!���C��F�0*R��Ɯ�T�ʇ�4��~�C��B"+[Yp9�xwB��Y��Xv�4(�J�0�G�G�!�bi�B�#��E�-���=�� F�������W&>�� �O�gG��Y�1���`�H�h��!I	g6H��H�e��by���2 ,��V��@*����?�d	�D�2�߱�@�$+�J�WطG�P�$+��1�,�J��N�ե�w���@��&Kw�x�$q���w_�ۅQ�D���j�
?�ŁP.��6���=�v7�5.���:�#���l��C
�ݠҩ���2[#���	]��L#�
G.�o��-jkF�o��^���PFGs���Z��>V�#T�Y�����p�Z��K&�-T���e��*l�H33�Fܡ���[��gU��)4E�g�ޛƒ�a��z5���/���9�Q�i_H�R5B-�O��K�pIJ���8�itߓ���o��~K�ٌ?ӀWS����gs4)xS[ \v�p�v�����2�6�Q�_~���H�R$,*QZ?J�\o��t��Wϋ�1�س
�a�H{0V�`�~�F�q�	��Q�w�e�<E��j(���7c��k�^}Am�L�3i�=v�ճ8�%Y	H��l�ڬM���H|,��b�nނ��7�� $��Q��H�QI:���&��y]{:��4?+��K?�����D���`�h���y��u���ʰ�X���R��0}��"�m���v:hrp�=<J���x�.j�p1\��wX'�:"l�k�2�%����S4j��=��+}�u&Τ�sL}Jv��r�����l�{CD�:��5���PXa�i�ǻwzq�W�����o׆D��짔�l��L�!��iԋ��1���kY<��������8������
�H�[eŗVx��[���#���2s�� !���(�4��^�h#+�M�{R���n8��Vn����C��&e�I��Gژے��AMuԋ"RBgn
lMG�m�p$>�J�g:�-lP�_OW"GV�����0ca"�FTi�'�nÔ~�0(5e��#A(Enߒw��EQ��NBi2R����8���>j�:����B��c�#���P�`E�K�dj���#N�`��]n�(=o��~���E�[��s�Ӽ0zl�Z@��v͍X��B�5�P���
��\�Qȯ���e��{r�-�`8�&p�5m,	n�.�4l�W��i�1R�9��c�@v1 ��:޿�H`����=	�g�+r�"�+����Bj�:Qdy(�Ǿs�G�1��Mei�Z���8a�H����bU6�Q�T�j��	��Y�zE���p��Í�u�jس� ��#j������,�ƒl�dfE*��r2>�,�~+T���$-[h�9-W�a�<�_� )Ɛ�X�b%� �f0U-������$�"]�(�f{�K��]CL��C%�Q(3I(�J �	{��r>q��jQ�Ğ4?���*ceezŃZD:O��-��6�0:��%�1[R�:0u]��`;v�h��C