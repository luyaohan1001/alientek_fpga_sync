��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�4#��71�Q�'���9�������uAg�'!eʓB�`1��_�#����(��ú�"�
i!酨#9 ���Y]�>8	p�  ���	$W�Ls��$�,�`����$	�p��[�S�ƄҠ#�yP�KuyD��+��S��4��0Z[]�i�|����
!�V5��"G�p�~��p����K�@g0�$��2����e �,��Ra�SH�c�(b'�Cό6r�"%�A6'��#6p�
h!�@��%������eV������c�߇�5�tF�8	��<z�[����x��JuZ�Z霼z�[x�mf�f����F#�BФ��?[g���#�:*��IXr�������ʇ���\I��( U��a�?�B ���.9�)�g0�G�����M2�÷�'jo����X�.�R�⻐����w��w�	��1����f㱜!ͳ �V�Ca�U�JB6.���8��U~�NҞ�>��l?�e;M~;�H4�?��[m 7w֋U7'g�V�&�� �W="|-���G����^��[C�_�{7�!3���Δ�y8��DYro$������w���y)�Gɸ�S�~��;x~Tt��X<Dw�Z�Ɂ&���	>l!bW>՘k�zmS�>,�H�D��=�a�R��0����M&3"��.��*z���S��?�L�kx���}��aC�R���{g^LKj7���w�us�	�`J�C;��C�R��Մ���.cǢ=���mn��W�'x`z=���Je�5jm�N���W����V��*�Ҡ���뢅�a��K}��X��Xi�2����ѩ=�v
xR�\��O��s���S���Q:��'V�����s��Y'Fj���b:��+���'�f9uJ��s�ۂtz<ng���3f_�j��z��s��G>�0\ʨ�j�3�#k�Y�ͮ�M~�.�E��X�C�R`/f���E�Gr���%2
��;�m�A�;�Of@/{5���H︕ M�5a��v���$���aef �i9,7�ĻKFT��j�����tԹ�s�K������n&�R�ȓϑ�pIX�31�4f�~����낱�[��$g*
>�T�ȤW��3�+ i�b~��3F�I�gAf �����ʀ�'%��0�J7�;9j2=6_��2�m!��g�nCQ�?Q�!
)�H��w�	ћT���+7��|�5�#��Ք�1�=r2��gR���F��jf/'���r��7�l��V�0u��eJs�Ȍ������^��U�	xow1��(�ej�ִ@Z���;5P�ڔ�4�U`��,���_ݼ�}L�W��A0r�)#�>����0]�� �J8n���Qw�7�j��j\��F��q��`�W�%b]Ƈgɛ���o�Q	V�+4��A\k��[�Y�'�l9�m�A���]�u�;މ\��!�`d'8o������uH��T�x��^DWn��:�TV2�E�o�LZ���V�LW�-�+HI�cκh8F"`��&a��{קr��3φ�Sڴ���� Uވ|�CYd�ȟ��G<��"[�7�����n�(���r`�*��O+�G�:E�E��K-�U�9vڎ�:���-�FJ�*�z���A��Y�x$�6�R}��~C4	�Z��C�ρl�⸖�]|e�f��m�E��F�(�'Kg|�`˥l�9�J�m�T�`!����#�|�}����M� I<8�J+�/��6A�ļ#��<b�T�Ly%�	9����k��h�0�K��L+�tz� YӢş-��%�O�V�5�J�H��(��6��c�����o?<f�/�h_󣿙�ڃD{���ExN��(A�`ױ`̚P���?J�`���%�-e�@ث��V�$�'���{n�9�"�xS:о~'k��҅$��L��T�"O��C��E����*��)�#�U~,x�|;w�?ٔBx@�F@T!$���'@�~�}�^��)6�\���T���o��yz[�����AIBŠ*��ٝ� �^~���GP�|�M&�8��v�
�����
#z�K\>n�->6�<�y/#K5����P���OSu�%���_y�	z�
T�,"@���J��d$N�pyMXK*a�����A�Snءw��_:���R�Y$O��?�k�����:�|]�Ό�L�F ��S�{�[�N�f\L8P�'�Rv��n`��zF�
��^t�j�H�=����7DkN����uK��4N��I@1�?
�̞J���[@H��=����"dW_�j���n8���vc���ߧ�\�������"�\��_�Ko�0�O3m������H�}�<9����X����h�#3���@ֆD8~?�C�|���E���F�j� �am��<�4n:�"�W����M˯��k�tZ�A�^q�-@b� �ղ�a��ST�#�'N?�j��jJ�S&�<+ŀ��1��{�tf�Gt�z��n�b亄����C��W�k�`!t���'����N}DH���QCC���V�Ex{w���F��d���CKGf#P]���KU>N���۳?�Q,�q�����$�E�F��P�����79,�1���19�mquu�aLN���g�,�Y-����V{"��JI:�0��`�2��M��:��@�nA����5Y�^;�W�~�@	�!P�G5-C�/X�Þ»����3Ũ>�991���#�����ٰ��_�\������N�(���5�rwWc��+�#˩�ø�@�Ve9ݜ��~�T�;���Jq�����Gb�J��rF�
���a�G��[:��%@�eE���A}�߿�YS sI�>J:�$���az���2#�R�3��y�:^釫	����L���CcO�O˓� �5 �4.�8�X~�/�2�k߿ �M�a��]� �uUo� Ue�����9��/+>LK�;�Mu����b{�
��7\ш���}����P�\f��=*RO������K��C9��EX��"��p$�w������O����9����3&���DS쐤��2O���a�i�L�i�@���amV�o�f��O�N�{�_�5�Bi�,*%H޷�9��oG���Æ�����R�RA�?W���)?��:��l*�i���2D3;C�'��s���7yC��i!=�Z�f��3蟇��Kr�蚇9���(��tL4ğ��c�i��ñ2�NQ�{�����彈ʆX��U�(�D~i��w����&Fq�1#�
��{sЌ�h��T~���l��;W��;�������y��$ʽ"lv���7q����&��=�`ߝ�������oZ��t�#�^�>� Kr����0$�jLG�( V�����L�&4�7���b��37`�@��bno��1�L������j\��![>a��7���;� L���w��i�s��l���D��To��%)����>IL�b�0�u^������u�YI��YuB� [���?���J����tb��K�P�ا�~�/�G���	�I=;P�������yM�a��z��vCr�T������kA_M[LFЯ��_�ȮhV�X	)���%�Q	<���%���|��kM���/�z�Cou�U)����X+!��n���2=�2r|�_kIa ����spl:�!�	4\n$����z1�OV��B,�K2w��c���J�ʶ/:���R��D�N�vȉ�v[��5�<B��a�y�����+�R����hNy^�����&���?.��+X;P���D����l�z��H/Eg�������U|yU�U��b�o�k�U[�����o��H.���o�{�U��4��g>ۛ�(1��zqz8��0B�0W)�g�3Z�	�TL����ݸ��;�4�����ctndN�}�bp7�ܮ���`�pV�*d��]�w�y�8{�`&j;[�6[���-�:f�(��-�4B�!�ж�2p��	���،��,�)L�v���ޓ��2 u?Lhk�f<$W��Yq/l��n�vB�P3�bk���֟�=���a�w-�=;�j?���3;�~�5�m�����h����q��zبʛT6ҫ����KLGA� ��4������^[�U~>�U��� �@L	Mf>z��{(I���)9A��~���D�л�X�x.Ss>ZdpP�u��w�3��`=�<�4����?n�U<u����+���A����n������1��܆��V����.�=�6�6�����M��a9��]��ֹ^d��?R�����aF��:2�Dp�;�/z^��O	�H{�Ч3�7]=x������cP+�as@A�A>�ZLqW�,��]�<�T�w�]�{F,���Qnݢ�AQ�t��	�5$��q�%z۶�u��-� &�|���,H�����jc8@�"�A���|�թ��Fge׃Do����׼����<��iF�>�}��ꉜ1}Jvr��вC�IP*Pq5��+�0�upQ�\�D���V�<.�G��9�8��{��VÄ5����2�*�Y�*l~'�z�LmBCv�K���k����To�� vzN1Ѩ�h��U��_)`�C4<��xI�ƬP�����S�hq�4���O�5�x�j���}/�]�h~8��K�8e|t�����4D�o]h�$�?M�*�V �:��9"�$"�jb�-c�ZE^J��- m��4���;�%����lV�DÛ�.�%c��4)�2+Ā�,���ᩭ~���;�wp %{\���X�@����W!�=�I�E\pF��N[�k��^r:��Ըt_b���x��'y5�.o��r���!t�-'h��c~����%�ܗ�P���5R��Y�B���N˚�JB�&O׍�Q�!U�Eʃ�fL�"���qd���C��@����89c\�ϧ7e{�M�M������<����zb)d� ��#0�f��4ҸP���ql���ݪ�٥�&�'A���-Pb8�T��H�>��^���Cr�9�O� .�_��VCH%r�WR�U�ac/����LP��ռ�=h�e��'����v�ZK��=P����| �~o�Q`!%�szN�v�z�e�]��HI%��L>hW��,���v�So>�+z�ִl����b�)�a��_[[�oZr��Qڤ�H{B������بn��v�u�POdn��P�����P�w�"TN�GC�Y�N��e`|�~i��}��WL(W�=���[�����͙Bc����nb��ڋ�^���y�/�N-���X�ՠ���D�s�vw�H�!�lo^iG��Z����u%n�	74�_"M�G�7�Ũ�����/�s�E"_�My]�|��o�������d��"o��?T㢈g��6�q���-��VX��%�|;�IL��ߛ6+'��8ALaͭdrֽ�t[�����mé}��]J�J.2ڍ�pk���Ҽ�d�t&�c�
�+�#��Z�:f�7=)���g�2g�F��]5�� U�	i��[U�޿Ňf�{d�� 8���Py�ó�-�G� �P9�R�Q<�9�1��>�g�Ьn���6D%W��`b�<d��#�,��u����ō��c֌ɇS�)�� �-��	j�p����j��aF�#�o�[��$9{���9�a0,���v���c�j%�4xs�$[1�E�C��XT��I��Q����m�2��6E�H��Zh@
�&����h���]������S���x�&��UL5�����c���ǫ�?���3m}!�����La�]�]�`u���K�����~ki����D��}?�$������3cqM�YE��w�,���!�
��J�i]�}�w�t_%UTh�l�/���ګ!I8�A9�a��:|
r�ŵ{*��qW��z�`,#���=�_C�=��AOA�=�0��;QHm�F�j������kb}(�����>�D:{?�͛gd���4]p�/rC����[�Y$�J� ����_|8��g!G�������0����-��讖��r�u�A�<Gb�MR��S*o��H���y��.Qh��k��Y����g\#�@d�2��7��	�Z_��G�3���*GA��t|���D"�Q���W��Y!F�vT��ĊS�ҩ�R��X27���z1ݮk}z>���#������7Č)�^c�dT������/�҃o�?�[�+$V۬zhٕp1�k�8˥���{S��M�eˊK�l��F���aK~��̑��������!�ع��q�\��^u�~T�բ8�v7W+�3&����Y���Ov���ypC4�#�����Q�QV�dʒR����V�gHc��(��tn?2�K0�W ��	�)s��M����#�ԓŷ�O���k9�Fn�[VX�~�[~��~}����)�C�(����*����M����j�����OMCm���v4y�	|�$��7�΍�s��?p���3jCS+�RE:��B�Ԕyh	1�o����F���	�oP#ft[`4S�JsQ�)�'�#�b/g&����EӪ�4�h������]�%p܇&�5�3dܦ�l&~�)��C߈m�(���?��\�i*�;�cL(�USC#QO�C����U��|-�M��`���m����"�Ϙ�
G��y���ö�4�곘=�|-������.Վ��yW��d�����3�MLיO?�g<�ɫn�κp3�]��}��b�1�e2i��->�Zak�KIt�M��Б���@��R�WQ5��.Ņ|ۅpKe[�������)�L����O>�|.��lX��f���7����xz�+pt���C Y���3x��X$V@�= ��Æ����k;�Ch~���I��a�l-�>"��ƫ����`���}W�����w���vo�a;{�su��J���4q�f�������������T��r`G��J@��S=z���,�j����4�db}�ɔ6 -�a��-�BX-����`�M�I��H�X���e,��.�_D^��%b7�q�^��o�!��მDvF��F ?��r�`��'������?�ڂr��;_���<:Sq�x���CzF�ܬ����ܨI1؋������xA�O���Fp�iH����`^,ؔ:w
-�{W�*f
&j�����P]$_Y�0}�C��8�N1�"kT�7�:�_<T�<6E���l�* 1���R;Hۓ+[���	����N�.����~^��껆r#� k���W�o�|�
�G"�9�ܕ}� ~�}l\������=�m�ǹUC��~�Q�
��s��N����E_�E��̐�W���=2Q֌�ܜ3i����v�r,�����1�ls{������g,;D�5��V��^Ve�
�x�SIy܍2��P)x�3�W�(Z�� ��\���g�)j]uYB̺[��Y�%�ot��<������̿�7�n�ȪY��+@9��]�TK;$�J����>*	;���@4*��������a��OA�Z��}X�֐�Js�5�r�5t6��X���x��_�n����;V�u[Z+׉��9�=���nat[���U."4�� ���������C@�XE����L����e�;�$�����k@ŏq�v��'t[>$�s9�ij4a,�-�-�iZ:a�Fw��Ծ>ׂ]��,�a�MC�_�P��%	�.�k�T�So�>\8�� �kDwx͗�#[�W�іZ�ev}8�=�=m�Zg��e���qO���:<���y?We�x��:��EB3�H/��h�8��a�*�_(7�3��xS�]֖<�<���7�bS���� �?pm��qy+��19�����؄A��U�hz���p�	��\��)B@�[R���A�b��g�!;�O$�pv�D�]�q�A�y�Ci�~������a��>R9w��9a�<N\�%���yw�x"�P�'��'~w�bT����p��0���!f���PT;�u<��c�H�#)�[�@-r!�@�4Q��������^�n�Ho��;��X�^�_����$F�2F�5����n��t��f��s�"'�+.����}�gZ�Uج0��[�m�X�q0Qhf�{��ħ�{��J����U�5��~��辷6ozFZ�9&VMv!W �W���
�A����_�M��c�MX�i��g��EvRj�/�&�Y�脒4�+�jbe=��A&�k35�늕 B�`���X�Q������W����E�я�yլ��R��$�@H*߀{�)_��2[ϴ4]�Y�Up����a8��|đ;���Z��p��B��x��M���"5�B6�D!IYˇ��@�B\*��2��ncT|,1=��a��`8j6�����&�����G-g���ʡ�r��J�Ja/��w[�e��CBd!x[xKtf�� �mHړM6]�~��ǉg#�~���<Hy��S�v�g�I�T�-��O]O[��[s9����,�� �#���3��;�wi��G��~3uq��=�`C�[Z��ʟg�Q�Z+..~<Yl�!�zIm���[)����G��0�k����ϭv1/��F�*����9�ַ��q����@ۺ��A��GP��B�����ǒ�1{��՘��!`ݖϮ�v����|5\Ǌ�s�&D�i=%e-�gݭs��_�2�����ʘ�z����XN{���" ��ڎ7-�4��+�����Z߂lX�7 F*�Nv?��t����m��7��Z�s�x�h�y�So:����l:r�X��@�Ozx�d��8�_K�S2� 6;-x_Xm���]XElS.�)���y��/�.a&0[��8!��#ڟ��K��t����E��$yD	�~��_t6#��u���6;R����'��w<���r]�hZ���߹��E4� �E��6v�{��
���I���w.��n;�ys~�$8�	.�� ��&��И3���&6Q�8I��d����*SQs�7�
� Se3��j��]F"�vKP5sTű�di⊢А#�Ќ)�`qF'�8+	�Vu}gD�1Y�X��:R��<�n�M�;������6V"~�D�w��n�;�ޗ8
��M*�/e�`��8���"�ٙ��P%@
� n�̝$�k}�:�2ށ��!����Ѥw�c��I����[���%僝������\�Ax��]���Z|�d� ���(�w(;��횀U��&LΈ�k�8}��kj>���+ڧ]'T����:�?�U2���+��y�i�U�O��g/�J�z,ҭ��ڮ��1[4��v�d���o��b���N��w<[�<�"����ԇ߰��*z�gߞ�؎���/Ej�c|`�0�0�X(&�u�i��:��e,�bDu��L��D@��ˠ�!ǁ&zP �G�f�b��F�����)�8�mx)�
�MR���-?�LH돞��\�H�ر�����l0q�Pj�D���'*��u�@Y|��� ۚ �}0�E�V����#-�aC���I���W�h�I���Q>����PX7o� �C����X�g5�N��r�_�m�^�����v�ʐ
�Do�Hg׵At�<u�y2Y"��p|"�^>�ޯp�GЅ�P�	��`@�p%N@W�t�/(UѭU/��.@� ��H|ά$uc(��NV�����jS��z�B�8����m6�Z`>��π�/-"����z�x�h(�rΠ�^9���ޚ��������My�?T�݄��muO�SSQF�w�t�b�1ᾚ����Xv�1�~W��&�E���Ȩ�|�M�lG�x��2�{�;����yB�'��6v�d���(<��!�����O�&a͡K�R���㟋�6U#$��b3E~�� 6�A�"DI6,7Û��S�i��\��ե?s�H=NS$6��8!�0��� �AL3i܈�Qd��{�G��K��9<!�2d	��dD D�<���N�/b5��߾�^��.�*#�T7�n/�[+i ܌\Ƈ��p��|Hm@3�����o���+�A�܋�'^���m����~��31��m��qpFYi�$��]�f�~(��D`L�1=/o
��⩲����8~8Q�w��1.=K3�?3@OV6�m����M�b _T U��X�痔�|��m\Lv�%M��V�vR���eɯ��#�i��h�����i튧����6��)���#\��J��3|�>�^L�|�	;60D�DJ��Bu@˝�2�P`��^�e�< ψd>����V0=���<���'5���h)��F��\�Q���ǃ
7�[�y�Ę�e/�Cͻ�K����X���C=�5Q�ߐ���s��u���ˏ�Y����p�,+�w2����1"�_��I�݌$��2ٽ�h�Z��9���"fB��ͻ5�W��9���>� ��O�s��FǇ���������{�k��WA�G�^�1�7��F���Lhv,hm��0������h��e�I�y�{���]��B`�`�bY�(Y��υ!�]���dX}c�G��~g-|bS����:qY��M%�P`�m�:O9�������j�7�n�ʻ<s)Jě@�=bZ�|0�y��R����Ϡ�x�����^�w��E��R!�E�k��]Lρ;)ġ���-}���U�σ����[��;s�v�{�do�ӣz��7_�'X3�U�'rtM��1���(ɩ���-�0�,i�AlW��'��T�6��(�z父A}�F��ߐ?��OR��10R�������/���_1o��;A�������E���R��#�ƴ��$����7A�5AHS�J;,�����'}v�I\.�鿗���P�&����q�+%xz*�Ӻr:�:��'ţM��F3)���6z�����Ǡ
�T��7XQ8�b�2�F�ҟ�����l8�t�G���%��\o���]E\`0!i�����Ĺ���jQ��{����|��!U�P��_[�H��j���w����<Ԧh�F2���`���&��@@,M�]E�I_�?���x�}�4�,�W��L�n�Pֲb2;�0s�~Q���!�~�� �	�1F`�t>GP��&X�'�>�X<�B���Na�\&a�w�X�s����%2��L�IBgNyMz�d�����S1[ۛ�\��;]��Ym�_}d;��M_�H�I��4ƝAXN�Z��Zӿ�f�MO�e�%�Y�3���Ӌd�i)���S}��(�`�7d�a}D֘+�PH�_��A&���ݣ�#�//��\�����$����a�A��:�0�l9���u����xC`�}v����d��dos�X2ħ� p�ixL�ҋ����E�V}���!��H.q��\X^'����w���
6c��k�g��"�.v��딷iq�{�:h���7Xla˂RV��v(�Ri̝/]�Q��*^�������v�*������?�H����H�G��6Q\
d%�NyR�񮹣0�c������1��g��<�������Բ�\ Qn�)SBݬ�FA:�ж��.��Ux�����"1t�&�H'	���L�Np��aE��zI����n�`�L+Q�.��{� ��Y �D�u���ݨ�W�\��2��^x�F�zDF�����
��lJ:����"e�������n: qHJ�|�R�W4���t� �c!�5�=�%���*�^i�%H>�:�;���ot��#�s����y��0�C��wԷ@�f7��~W�g�����JƔ���@;@vz��\�֚�2�],�Wo�gyD[�6h��+��־m^Pp�I Q�(6;��+{�㻒{�:�i��v�{��&�VH \�7�����EN�~Q�|m��]�K�C`�x(�pF���Yf ��Q��_@{�xv�Ҝ,���nB���e����32���%����G ���G�t�5M_tI*Α�	~g/I5D�f���T��-4u�]'3�z
���Վ�w53v���v1�G�����O���dKH�	���^�leCj�-,'�u#6J=���S�K��UfK(���w�1j�0`��s�Ki�����s)��o���_��^�JV��Ѯ(�d=����;o�M��0�j��
�ۆK/�;eD�����Vj	'� �jO� ��W�(Ԅ�S��=��g�rvZmH���I ���pB}U������L�(��>�V�#����Dh��{IC��Z�ӈ*��2� f�~��0�n�l@/"k{x��e�f�.�����E��m:�`��4�/Y�P,8s*	mx����ѝ.��r$PT���=L��ud�g�l���e�6���҄Vo�s���h8�������m����S�Iݤ����rD���m��au�����+�M\�ڇ�փKHIaM�B��E�Ԍ��J+$�/	/�����{c�Ԁ��Bg����c��"�1�0U'*bk�v��������Bb�(�R���Rz70��ʁ�&��� �s�s���f��:d=�W���\�Uʛ���3����+,Y�_T�8��8%���ߢ5��$&]�z�ԗZ��Q߁>�'��'�J�4*r��<`�11*g�T�v'�F�S�0�R��F�b�b,wZ�W� ��ɮ#����h���r�����������n�R:��x��n�姾�<6RNG�Eֹ%u|��5�����Ŋ���6�P�Nb��H9�H�!�� ԲC��r��9�:�.�#�R�'6.G0�}�!&H53[Wecqb�mvi+����/�]����`��/U�$�M<L��_��L������wuL�2��
��׆�"�wny���msQ����s��d�5�����?��C���}���I��$�܇n�<�gM77oZ�A�+&F$���*��d;[�u~�O��`�O/ga���2�P���	��iF���*��p�/CX��w> ���#�[�TA���ݎj��Z�&$�͢"}����@���C^�X��~���c�����ޟ��v�7i�ƐZ���ď���B�P�����ᕩ�����B��c��Ni�w�������]�}��Ǻ�N�|ˮ��T�JQ�3���\)�ƚ7�=�%�	�W9n�k��Y�?'{��"'�C�/�4h��d	y�̟�hp_|�v/�b�(zd�y�`���JC����Mj���α��l�z_�,͈Sz<}I��JC@ّΩ�c��y"Xp��:�[}Ql	GI���
���ҁ���XQU���0�Ԣ������H銺^R:�����`?8֫ʘh��@Y֡���t�����$�\1bfz����:CZK���l����vcޯ��C�e ���<6ipO�pTJ5\��CE	n�5:���Ο@��Ԁ�@�/TC�bo�w�����BM땊�+�����u�P��^4Q��(*�]�4<zn>�ؽA�ZT�+��B
�b��΁�@C�@�n�&$��0�TC/���+��q#�w �p�v /���Kz��5��9�^焷�c�
�Y�E�������$z�l���Q��o+�
��6u�R'#X���\q�\�&T(�q�P��ģ@�'1�͗D;8r����bl2�d(q�����,ɝ�ڂI�PjN'��px�34o�����2�W�s��#áC�x�}{L��D�:)��ި��5�����lW�2��VN�������G�o���X���j~���h{��ʾ�{bV�*	�!��%���l��;ߕ�(^7MG	T�?���\{�4�#5!�r�av����51:�Mr���m���~U�`@k�ѯ:���3��r�~>Е�%HQ��<����KMCK
 ���s��G��.�{��+�D�����r(�'i��'m7�~��!v���)L��'��|�:\ ����:����i�q�QLf.#��'`���2�-1G�;�peʒ���19�J\�y��@�O~��*b\�� ѣ!{͋�����������B�2���(��<��o��t52�Tz�a��A����|��F�	x��؄G����R=���U~ʞE<E�d��z�a��$Λ�6܋Z6�����(3�h����\EU�Iq�����3����Oٗ0/��W� ճ=������h�m�Nύ���qS�@�Zעj��!)�B#E�G�8�����.(ipـ����a%v����/p��x�)R��n���R6�]9�n`i������P1��a�6��K=�ulӑ��R����Gva��/+Wώq#y��yFM�"�ʩξt�fv��,�����r���c����v�?v�z*��q:�h�A�HG���	N%̶�C��>_ �'o�onH�*>�`�\"r	������Eȑ�޿d`��ֳ茡��f�G�K�����ԐEB���I�SW�i�as�)��Y�����=uGQ�E"�'����_Fu/@W�s�2�G�<s�aq�Xp����(��H'��ߩ��~!��>+�A���jl�k�F����&��0e��fW��eNm��N��c~�5�!)�m���'�,�.U��,}���T�FE�
ʉu��MWI��/ݭv>zV�ʆ���04�gU�?��b��ޔ$`�B��k�E��Vhg��uU%��8�e^^�����8>B:&�F���i��us��u��֕�$��4���]����&~���Q��`a|]L��7ד��TQ�t�!i���*�9�z
Ӛ�ݛn�os�F�l-����#��F��nz�S�y���^ң���枎����9͌������I�L��Ta*y�Į�P���߳}Ֆ憅d�s���.)p���V���+�*�;� \T5�t�:L���2!<��k#y�!"e['^H���ch��Ch���7(�7Vۓ��%�KE�f5<މ��{�4xBWym�*ن��O�_񤕰҂�l��v� �[��q�)?J�K��*������Ɔ�D{���$�l��d'H��:�E�ۋ0����?M	y�Ĭʞ�se��\�{��%{�'��^}�B�����>e�rzohm����}/�j�븓o��C/R��LP�Y��-$/�W��	��9(,i`�T�V��D�B�c�>��ތm[&5d��pP����O����/K�Q�x~W�ʉ2�5�ň�N�������c�ǊD��� ��g0��nn� �����96�l���Q�@l�ʰ2��b�AB6��'b$�.vM��Z�'HX�Bk��xP\X�.�!<Z��ր����b�$>[����4?�ĝ�P�W�@�ް҈��]
�}j�%�����`���-5���{���髂s�>(oÀPT��<M��BT�+��X�6�Z�4x�rNq�^!1/y]Z�u�ڨ�+�lͯ�Ʃq��st����:����@\�-����`��A�?�B�q籉p���V�wv�@��ʂ��А����tL�\VH��͢s�zT��G�LG" �q���f��EȻq7�%�
��(�.i?��U��a���C�=Ye�ei�F����V�d����H�x�6�#���}x��!ED��ӟ�v�f��<DG�餫Jx%�<�D%��sy�ρ��^Iz7 =e�W~x���g�W�T݅�ػ���h<�8�����˻�Szf�������k&̮m�=cL�Aܠ�����&�� �YA��������XBՐ:Iu�"a��6�l��&_�I�g@���Z��� ��,�{*��0���ضA��$:8�/�o��4XQJ���c��������ܵ�n�\�Z���K0e�M�B�nr$���]��2�sϴY۴��I���(�
�Wj�OMD!���8�V�:p�lM2�����R�w�5m��
!��U�+}L9wi��]�qZ;Ÿ~��N<���0q]^<D�'�ȣǮ'6n����k�}H���W�ߐfV�����w�d*��Y��RfGz �����`��s#����H�.���Xݕ9ѣ�c��O�����{��c\��n�s�N�.	�9�1��t�t��i��?�H�|�}�E�S���tcW�ژ;�ɏ&��nZJ�^�ه��l�+*�O� Xi�Ȓ��i-5�K����v���������(�!�N��:I7��¡K��zp��'m��ڈf�@�Lp�|kQ0��o�	�I���Ӷ�����}��f�Q�f��	Yz}M�Û��IӠjG_L��,��
7"N�N�2�>CU�'���9�����������_������l�����o��KD�qol��d��Y�嶻 tab�8z�Թ��r�����_� ��6�3��U�7^��!|����'_�����1�<u�Ԥ��h�B�\%��;�6f�aa��֊�;�� ��_����kn{U@u�W�ӂ1�ԩrga�=��Bd',@���u:��}~o@Կ ;-o��>1��+	d&[��}i���r}ް�;�Y+Թ�a6��Fn �׆l�L,�(��)%?��X����vq���w���Y�fꪼߘ�F�Z	VnEtb��:+K�gF�_q�X�A�:b�{9�	�)>
��4�����<B&�vP���0�@�"=�Pf�&Uq�m���)xOI�jS�������*LxZ���wܩr�[�Q�y�sG_ҵj�����
�_����ވ��1[,�nq���r��rݶ9�`:t����4Qf'��{�Ơo�o�`Ft�/�^�h}�Bd����H�>5����<*�Q_82����(#��s�C�b���j�r��b/&>C��0��������܇�7p��ş�j���d�|�rs*���i�G ��t��y*1W��<[��[�����Z�)���AX����(��0�g�y�;��^����+\%���3_��h��w��	������H�8��g�J��~�d˂�uez&��W9'([�,�D/�_3.i��V7њ�#���I�CU��p�C��;yWsڰ��vR�Q�߰��f��L�;J�s
p�0��N�23i��b׎��P��|�3�N
�0ϝ&?B��ܠǀ$�m�-fI&��̼��ZF)fez�O����Ū�nƯ7](���ȶ �u��� �V #��	XxmS�ecs2��XrE�ͱ���e0�ԴD,�8�c���F|[%�i\	����Uiy���=e�\����qO7�5�wza��Q�u�7�|?tC�@v����k'x�et�����SGn�?����_p���L@�8�)���������}&���p�� ��	��I�����{�C_��~���(JF�ges��d�����N�>d�����T�z6a�[x�l�1���08��l�ݨ�����}��uL�l���#��%�~K\�k�
�E�Į�H8��e�׼�<x_=%_fN�Է���fQ��������t����'z���BьC�Y�@��o�.��b�: �mmz��A�D[!�NHyp�'*�'BX����j�T����|�î>%04�5z���'��9�����Jw��T��E���e�	yrU�g����M�d
��ڕT�b��3D�;�?�������r�?��ON&'�eB�p��!�o�<{.o�����d����ꐚ����E�6L�?�:e&n���J4�ͅ�5��R���}+�zA��d�� ���!��j([㛒�8"�y��E?�P0eM�eRx�z�
�|���<�eQ���Ɯ��A� ����J��p�R5�0B��vx3P-���;���y�kI���v'eƢx@g1xy����m_�Jp�dc(3�e_���`�c�=x�3½���}+�s��$.HQl��9��f�����JO����LT��T�/�o�. .�[���:�B!̍�>�e��W�Y���5�<��D$�}����������G�[}V�p+��H�5����L[r�Lo�#�v�F��{p����ٟ�aS�Fr�"/GPp�f�m#��WĤ�������xRj�x!WjL�8QzZ�hT7hF�Z�m(%K�%����p�v�\i0�N��zrU�6.f�8XP�)^�]T�)CG,�\�s��I������Q������	�¢�c/�dߠ�9�D�>#^ΫR��T��}�C��?;�}��8��₽�zeâ6�$5sV���t�؎�� ��)��l�D�!-JP�KH�'��rn�nIz�:�>�!�b�����������"ogi,�����Du���{F �V�Z���;�%�oϑ���� ���J�;���(M���w�9;�PG�Ug@�eظ�����L���O��2���K�]�*R��e����t9�c����q[�b/bK�����I�Mj�c1>��Wfd��&j��r�*�P�c���Q��~M���ʬ<�3�%��X�q�l9QeIi�E���sOQN�t��{��WԎoq
�np��͈Ŵ���ɢU Rd��2g�2�d�Zlw�k�s��R�&8l��[�H�@�^?�4$,�Vc��ɏv>xt�'�������0�6p��&�R�u���G�wYG��aL>��廗�H�T"�r뉁�6e��Wc
�F!a��~0t:�<�+hH�z�9N��.W�ڳ��g��{���ޖ��v~>]2��_��x�j���n�Zy�m�����k�t��ezV�-�Z�S�ϓ�RM�5A�8��.�Gj.�6���9, )����)��߻<��a_Vj�J{��L9��++(@�,A��Z�:2���j1F�"�K�9��{|l'�����+b�rn�S�������[���_�>:fzq<�X>�G�1)3������~S2�B�wCU>g�d���3,�|
\�N>�3w���\�JT�דԞ��r^<��Z�t#�#���z:�㇬"�0�!�y3I�	��-��z]�c'�����D�E�◌_�u�y���,ǿ����0�J��+��1���o�l�-D���Co25�e��V ]�x�0{�T�<��s~<$K��m�n����c��@y^b�Rr�2;ʎM�y$;O�=�
C�����f���U!��=u�H�V+r=N]+���E�-V�n ��Ef����G-�К�}dw���D����*�����2���~��I_��\4�L���5��"�eԡʻ��9!Ep1} ��v�&Wo�6©G�0��H���M>���7Y�r��":�e���"Ɩ�Lv�8�e���������S�(OtgH��~�x����&uS�*�zUPX���*\#����\�S�s �h����dY�1%1�]o�	)~�E�1��0޼J/�aH�9�y���&gƳ�s����>�<�����|�����²!2�]� 7�td����BZ�O���q���F��=���,�Tc/ZN��ߺK?�+'�����L�T�4e��Ѯ����z��chu "��L �=�	5I���[�K�tz�=�cw�	�Y�C�!�+S�0�N���,��ޭݒ����*�J�v RX7�&�vK�E���Wd���:��\.j!|��;Q�Q�t4�Q�ҭ�S�YD��u�}��D�ႌ]?]୥�QP�\���R��C�r���'��Y�NOӆK���^Ͷ��*C6p�.�ϛ��x4!�[H�<��NK�_Z�mH+����='(;�T����J�3_7����xc�;j~L3;jWm�� �)gr��R�״o��kƃ��E0Ձ��MMm�������Y	Ѯ�u�7y�f1r]�8�H(iXo�w �o�?{��s�2�f�PI�B����w/=�̼ɽl��3�R�us1#C	� {E�D3�-�B����jZ{�mrR&/�����(t�FV�{���
=o�@:�	�������@��Ȭ��l�٧�<~V�(Z��[E�T�m?}�d�-v(4Lr��ti����J�.� �%�>��I��-���*�d���ʤ�Xs:��X��G��K�t�F#�"上}��;�
�<����EL2ݎ�mQ��\U���Nb��c?�9�v�4�����5��
#\sNBq^��i�ɣ!Fϔ�"�~j-hG��K������H;Șc��=L�AD�}�1%��X�H���?.N��z���Tb�v�BI?A���EkH;H�+� �*Z.'GT�9��U�#5e(��_~۞^�����N�@_�����-k�*8�7v�v�T�e�_ioe�P �
h��ƫe�0ω��NJ$����4��o�C�Q(�Y�פ_@e@���#����PBTX�hm�Fͣ�"�Ҏ���vdW�G�O0VB�{(��+'�4�_�G�/;�#zl�ST����{�0:�z�?�f���Q��.09�GMT�T���:��o�}����F1(���b� �ZzQ�M5l��᫾3r�]]J��)�ܾ&ٷr{�;�E��2�E:C�iy6���'!YTd)^)��x�P���tb˦��6a����`E��V���g���'56�۱IZoE<�EV����*�B�O��M�1���u���ϒ��~D����U;�!�U�n��7\��9��2�$ݒ�P��jTT���9���� ��K�d:�w:�u�(����������-�� ��3����}M�����.����}'�!LF�4l���4��#\��/� F�GB��_� ��<b[֔��c�%����N���^����3q �<����:s��ډ(�=��v�X�Z����0c�f�
n:,z��(4��-�}�s4骬/�a���A�i�=  v���ct��t'�eic�քD�E���̲�K�Ns$\ϯ���"�;r�޻�C�V�� (v��֬�3F���d����?��ٙ�d���<ɂ����$/��A�
�_�v��T�%^R�Q�:�[�m���v.Vkn��L�B8%Y��Z2�{썢�fؒ?��QU����2M����-VQ;����c�0A��vBZ ������#*�j��r_x�`���T���"D|�;�ۦ�Ft��mC/I.�i�i�"Kl��d,�o��?��w1�WO���x�� 8�n̡�g�pE.'O�9V	C��G����7�6Je{Չy�/�����0��RC�䥯sǭ�bl������S�,bG�4�?s���6��/5�홠#��U]f���N���;BBЎ�'��~n8b���f.���r̦(і�,Ie�zV��<R�!9��f�r5(��~C�R�mX���l�r`t��?p��%�]!9��Ǹ���@i4�5~����:a����]*%&�:2�]'6��esO��#H�P�vTk�x_Ic��"Tx� ���-��}�1�D)>��Ou!��|�$Ix��T�@R�.X��zy��<�x��x�E�.vn0=	����y���J$��y{��.Y��g��xZ`x�xK/fd�D��;jUa����v��f�䌫1����DZ)��ؑh�>�N=5*� �s��1�=onSv��*O4�t�M�(�+d�f��6���g�k��o�P��&��wц��L,��;��R���U����J��i�Co�2�@ն�>�����k]%,�8m�� ��#��t20���#yii�r�VԋB�.�Җ�o'���j�i\�j�������8�
d�vW7Vg#�ÝTb��P��"���^�~j�7��zPWw��,�.-��<?�d��t?��3���P�F�kz����ٛ]$@tJn��F�8Nȍ'�˘ȳ�I�!�%����ؗ��*��+��j/�?��9�`��(������Z�%��������83�&=�41�WĹINI��Pͨ<�줅�o�����{ni4�`K&�-�+'eF�0�<�������Ɉ²a1���c6��P��+��kH8c�\�0w�K@8>|.��'�&��ܯ�,��!���5�=J�����^ro�JԥB�#�:��'ʥI'!zsh�im��JlsZJ^W��k��z�Q�	����;S�;
�ʧ�0�	�kI�*eM!�y$�_.w����s]�����_5-�ܷ[��d�1<0�Sͺ�F��N�lN4F�*�#߀;�RLГA��� �H�K�P2�mJt�l��Á>"��l��|���d��<$��@����*
;8�"(���0V�O�fA�g�<��'i����$�f>��m)y_�?0����=��Z�t��y������4��%gNRp���5tO!Špu�f��$}����4(���q���2��!M�O�S),CT#��*���|�.gYz��$g� ����=���(9�M�J�ȫ�җ�6��u�\�z�a�/���'��ܲ�*���0Pg�G:�F��m�۞_M���1�0�ŵJI�&8��'�OI4$G'O�U���rf�=B�{�~��`��]�
�[��� �ˀ��0�<!'��M�80T�b��������������	� ')U
�3�ʕ$ӵ츇뎕���B'c�b"�0+�Y6���*k��eh�{��B��F����� ����X�&��K����!�[�P��vE�l��^�!�x �lx�X���{1���98h��� �,�7m:��/��
QOz�N�ڀﲸ"T+(TC�K�q4 �_� ZċM0���l�c�޼qj&�+�� ��1�&���d�']�U͚@�3X�����~��ׁ���t��p����bG�Mn�Ru~Mc0-�f�^���9�f�|��:����n}B'�%�}Z��F����9�+zZ�\�%9>z�!�T�&x|-m��F�@�Ҋ,/��\�&�[?����/{�t������hv����C���N�Ivh��O1������Jۥ�����r���k��^����}2�s�F�!�z���ӢdA�!��w]�*E��Rq�FRv����&#�k��'V'�p�QVk6����ܚQ�ք�ڵsx�~��R��4��,�}O�.M�~�/���'g<UwKS�@���,޸�HU�R�a!*����>}�j�� Y����&��r*�X�#�C�Fɏy��o�z��k�b=7�[h<c���!$�f��M��Y���.
�m��H����k���C*�9���h�eΩ	��fi��	�h215����E�q;i�b�S{�8̨퀯���3��K=���D@���ݍ���ʄYMΛ��k�3Y ��i�z��K���h ��ޫ��*��AiU/7&�*���mm�p�>�D
�B�n�|$p)�D�]p�»4UR<|c���Hf�����{���"C�}蔙P_��,�( ��≭3ɲV5�I�^���j�q-���j!$G��^��&w�9p�q�o���m)�Vm�z$Td܈��	�>0qV�^9�4�e���e�v��y	�����6yc����X��,?R'���ʵVJے�^ۗˁ�HG���r�(\����6�bb�r�D��(ǂ�1�淽�Ï���k��_�x�#�8���*Ń� �44S�g�p�:;�g��.?#�Y�?���
��D&��qO]x*�ve��g&XA���)���*0��W�v:��s�j�+8��݋Cc�-�;�}q��eX�V�}��*�Z;bm�)%O(���4NWS��� t~K�g�}�=�3Ȝ!Y�b�E�
4�KAˑ����L�q������͘4;�l'1�׶�4�,��XI��مp#h���n������qhQ_�l$gj.�O)���tAN5�ٽ���Eh�o��9h[|T�`����kzǛ�5�p�	+i璲�
�#)M��A�ן�/ �R=��m���Ø}+�T���Ӽ�{�7T�&S�}�䀒�$������x�����MJ�"y�|��E\�g�\;�!kAb16팪eY�:O�96�j�X��?�yBe1>{�J�5�$�l��[��,6]��d���t�Gf*������A�����	v_�ѳo4�h��N��E��Ų���[��|6f���x�mC�:|V�\Ve�Y�T��dyz6��M����6t�R'�#� <���xv� ���وg�N��"�v�M;U�Y��p�%���>?�>OC� s��4�%��iv_��P�D�AS�xtK%�~�A�J�v�=n0��/���� ��K�c2����q��c��14�� ׄ%
�x5OG�w#?�grvA�h�ifZ�I�]1�p��)a��ȑ��(X'���a!ܷ?.��
=㹯�6�����[�O��8�_�:��N���%�����U0��u5.�ߧ~]E�e�&݁�$�gU��a�� ),կ~���<j�:o�}v�W������m�#?��u���.q�����hD�*u�r~��������G�x�̈́���f�l���ۗ���4��=kP$u�@�~��>b%���dc�FY���~�a�O�J�#Ye�����E3�
>�� ��L%�g�Znv�@��<��s�n10��7�^���-F9�yq>9������!m�����)R��3B�ǈ��LF��z?�z��<����Cv�`8E�/�T	k���b�b��7�Z���C��U(j��>�.X0�/����f7@$X5�"QYnP���J�x|u��j�����o��7mg��/��{5�;�|�ň�p���Yv�ܚ�Z�3A0u*P71|�d�?+�S@lߝ;?]�fĲ0���fEyw�s��B�]�C�(U$��)c�Ji�QqD�W)�� ״R)�j�����M#�$���L0V����j���"�k*�'����Ԡ3� �l6��ْ�����]���t����0�h�Ev։ଞ�3j�},7����k����;��N���~�dph��k��VO[e��Gq�j�Ɋ(+ �^��.�Z6��G�:��=�t\1��S����1vڅ"�	�:��*��?� 8�2hyY�f�ц��fMd��r����}|�M�N2��s�u���
j�8�r�0�H��� ���Y���,���e7|�N�-��`;���@	.��13�y5�����e�J�����w�@q��"9�E���]�,P����E���_xA��&�D�OZ�cd�J	����6�~ ��w���G���G8?٢(l0F�5�5ڔ󬰏6����&N����@<������}�H� �A>Pw��b��Ye��4ūăb�{dehi��mb^���dT�'^Q6�oz��bFeS��xi}��������kv���\_3F5<�x8�	l01�����W����p�<�+G�5�Ye�bo�|�b� �r=J �ou�a�]t'F,^��Y�V�n���z_��̥w#ER#	���_��e�V��ԣ��dB]�`=��w�qwl_�o=���-,fLW#���g�=���u��o1,�@�s��hPu�FS-(CD!�DL�B:����V#�nm���E���@J�6 mY���jy��ќ-�/N�+�袗�ST�y�yؤ=��P+_�Ϗ�̭�c��˛Ko^�.��%3z$����9�����?��е� }���v`XʓzFR ��6�=��r��$x,�ba�l�O},��D�HW4!� ��C�lְ��dS�dM��� �M�즍���?�*7 C��}q��b��t���w ��K��Kr\Yt�v�8v�2�2��aq0�ԍ����#���M�6�m�Q�[�m����d������[ɯ�4g�����.�$?����r�ah.W��@��`�*�r�	qW�D_��"��A��9+f>���Q�}�� :�c�y��*��.��KC�/�!��[��1�Cx��b9�Z�^�`q��f��>+����:�o��;�ΏZa�}�;Wp`/At�4�Z�N�6榗�u
9ȡ���BԠ�Hv�S�ߝ����*Ҋ�K�Ĥa��d��c%ӊG��H�I�e5$�lu��.�u)|H̆�/�Q�ϪNO�T�/?�o`+g&�ii��$~��s�d�Wi��ć�������l�dP�m�=����+�Ll@iU	��9d��5!�z���nT��SD�R���8X�I����}#���Y�I��R��I�v>䠧
yY
~wA����磯袢
�V�u��lTS��vX>�		S��ھ?��Ri�E{էC��dXێ�m����|n4�^��)&]�hP����eƁfrge�����ь��=l����l�YAm~������ay�~�!�b�tGn�n���qu7`g/V��l-���ԼI	=�&�m8Y�3�`�I�r4�e���.w��k�b)�ʴw�L��I�������NU�����Ł�i���*j	⪱#|�\xs87;p/�\b�By�9�s���;C���/�F�J��4�"�;��o�¹��z��2����e%���,���h(�V����^�2;�h���<
��P52>�V�����>����B-M�����t�������C�{�w��!��V�zkj��-�po9�K������Z/5�o�L���j��?\f�{A} ���Ǟ��/[l�p��h�u�P�������y%q�$��I|���^L`��
F������:����h���Rk����x(M���w\E� U����p*���s�Ip�v!�!�*7ϐ��c�؈z'��u"xd�Ua,�9�����$�6�1W@���;���
�P�qd�0�z��Z��D�CD$���+��B8b(#�z�i��E��W֒�[)f4�������&"���;F�^�^E�4��(���m={h�g�B���?�bn�+Bd:���49�}�i1��
�}�G�(���H�#ޯ����¾o���k��Ѣ����"���,���I�`'sux1��:=-hy��z���owz�Q��̂5Un:
R���\�XȢ/�^�u���|�ɽ�{Q�H�G	7.S��LIY9(ֹ���md>�����(~��bm��ڿ�*���v+�Ի���mhlw)z{d���B<����LS|l�(H�t�u��D�HC��� �5xГ�ˮ�留�&Kǔ���}�˽�I���΅̛�#�-��cN�4�b2[�р�`��;���E-bΖ��I��h֦���԰'� ���JG��<~m�e�MW\�R8h�!��P���C=<Sp([�==JB�+�W>�E5K�o�2�7��> ����@,5�!:E��9�v��	kʖ���2��*��	��ۋ_��iGv����f]��G��g�J~H�o�?"�/)�^�ñ>W����%BF{8^�Ly�W).�/#%��e��b���=,�o�ݛ��r`!`1�{-_�p�?��]f�(GU�R)&�F&ћ�����Ĉ�5�$Py>u07�dkj14� ��� k+�r�a��,�A��Ry=�kɕ[��m��Lx��dF-�d"B�a�ipJ5�>��g:�˂sDh����)�E�/^N�Ú����}{+e<;F>���XD�.�����F�?ؐ� �C�?!eO^�+�҂��d��	�M�>e��%D�W�0h�%/�mՒ�]���-L>|���^��NkQ26���t���!����*@�C)O�g�M��Pȶ��*�X{c�)�ɻ^-��9ݡ�ց�rܳ�f`�~��C����eQH[��j�G7�b�r�
J_����˴�[�~Ж�h��ׄ:� ��Ǧ���M Q�qo�f�@�;��;�m(��oD��x����f6�Y�ҍ��fX�k4���R�d��1�2���1�y�)��|em[.n�L��]ZZ	�����lV���?��N�&ԞB J�_)�<��e�Ra���+��^P� !te����)� ,MD�M��#&�p	��7�Z%�Cuޒ� hH@,r-�����}CΉ�~�^L�d��ئD���gΫ#yLb�Ht�,�b��q�uM)񙫑0�jX�Q���@R���L���[�xQ�C�KR_�<����뉽�
V��8��f�֜H�o".�J(&@U����?d��&�R��)�n��7����8
����TΔ.�����]aV�6h�z����+��<]�g�#i�1�j��^�y�CְT��U��w���Cyҝ6@�y'8J��Kj�hn���FK��1+Jz�R�Zq.H/yu�"���/��G����r��Y�����H>j�,��0�?՚q�!@-@������ɣ�D�3�#RN}��6|̹}��D�T�=�3	E	u��j�{����lT�T��+sv#���d�Tu�r��tg�V�S3�48I�ݨ]���Aϭݜ�n��ɝ\˕���/3���EX+	9>�����%�������e�Y��Z�����_K���
�eg��į��v*�
��~�Xr������3��
������J��*F��+���ߠD��E������q崛G�<�����x:�6�Sy%y�1�y�G�9��Հ�J����G��O��i�MC[�`w��z�g���p&����~*��M�8��C��T�|��َ�����K�s���4z�����w%�UHfr��5��tI�
q�\8�C2����cT�t\`) ��
�]�������-o���ܙw���?7�ʲ"��7Z#t����B܌-���hv��ß&,q�^���O����ES�0����J�Y�_�(e� ����tK!�O�~��&!���4�d�v��+V�7V�F�Ѭ�#����x�%�d�j�;� r��[*y��ZN�%��O�Z*�8�vn�M�b���{�<=�'-��G��V�}� �grh~�t�k}�I1$,��bau������H�!�܊��� �zP1�A�I�o��v��0�93�?�E��z�>�H�G�@]��S��	<Swܣ��pM�|J�#p��������&�@ݎ �? d��ԟ,����	cNf��%�k�!3���@���n��z|��s�yʛ�~mH�ߢ`?Sv�;�ޫ����L��OϿu���]ƭ�BT� ̰�n�1�>�D�,��i��@�_��ە;�m�����=�<�_C�IG��1C'��k,���^ۘ�_���'��{����@
'ƓAE�ϴ����z���N�p���Dᢐ�O�^�:y]-FR�	�>��-��[	�h����p�M��D���5�`���86l�|uc�ܒ�E����=A)9C`I�iTe玣�U��WI�#S��{b���0<\P4z�L&�ˢ�D�㬂�a<�v+.ﲸ�\k ?6ϵ;�&��9�#����x"���mx�f�B�w��}�����g����Hv�!T���gKOX��Z�u����p�r�Ƹ\9�B�?ڧ�u;پ��Ĕ����x�.�Q}h��ؘD䍤���$x�*f��=��F���r��Uպ�L^�h�̦��8%�ә�	_sf��T���m�i����{������O����pIr%$�C���̸���E+c��OV^·�t���B#v~y�4��������a:WZ��gj6���<k����{�l��s��E&�zV�#(suh��w�gkg`����Ieޤ�*]n0	U:Z9�R_���%*k'/�h�[,ʺ.�t-x,Dv�OX?>�We�7D���pu��;��np��G���2���Lb�FJ�!Rա5�U�I�_��$�?�{���Xڜ�L(��h���rG��P��k���W,:�=�A�N-�6�!�qN,���v#U1*ęc�}*��	g�#l�[`�����~kX̐/�&AJ�\���?BU@[�w|��BK��̶_�S�2#C��1�L�R��Q��ȵ�������獐:귀�����u�?������d85�i���y�O��.��E-C��U�r`3{�&�������Ҕ8�$�����p�i�z�D���QP8� �S"���5N]i"���O3OCGN%�kd�+�țԔ����$l%�������<����4������o���;�A!�v$��4�W~בP�.[G,� Aǿ�HP�bXn��Z0�@4��JmpAG�,��$���h��<�z5��nII��|���;a��ɝ�ؘ��䡻z�q"��l����������!��:�	�}�lh'��w����rݶk���}"�ެL�^�/p�N�s�m'�q��<� g���A�d a��B���3"����-���2��Ӆ�u��婄����©�2[�3=��u�}�z��:�"
D+�'��(c-�gS��ξNj;ej��Ό0FT�e�o��� ή��Ycv�����X����@���5]�����]W�c��T�Ϋ%���!aq��e�ʴ�]x�\�X�����svY�M��$�3P�Zy�O��>Z��������?���%F�Ej�F�� �G���x1�e����Q��ӛ
����Bm�G�1��Ώ�!c���D���G����f[V>�I_�T �,�^*h�g���R�C��^i�|c\�Яd� �`�.���-7d,d�yK$�OW?5S�hn)�����<�m���חE��b/��<��Ť�-*�<'��:��w��w?~����gR�1�Ʒ�ߎu鱷�խ���t��Q�������	=���@iE�KJKX�Ӵ�Q�2MAҘ����ܰ���${�ND��|YK��o����,>�`ߪ��ϔ�ԣ�<���c�_����b�1�OZħV�	�}�H�@�9�Z�W�����v�� �%<�C�ܼ۬��'_a�t+�*��8�����p(��'F�p��-� `3��f�zd�������(me����%�(G�������h��MS����J�PN>g����y]t~p@���җM`4��w`�K92���R��1MaT:�zI��0�=��y
L$k���~�w�?�j��>�L{%{v�3͹Ԓ������mm�HS��b
�f@�܀{`���Y�������gk�G(҂["�?%�w:���%�c(����m rH'�Y�������߄55���v�b^G񘨌�?*(�����J��o�5qA���pX֞���H���,7��i,Y�I���}�/������yy\��}��y��$����L���-��-j��Q2���H��Z
D^g�B�g��n��&��?�m��x������dK��zW	������!��p�l�E�`k�L\w0�AH��X(��uء�����ұK�8���=WI�^��d� ��u,c�<��
���&��6,zk�e:8R���a���{zN���8��K`O�~i����S��R��Kr�S|!"ލm#�r�p�H�b؉����5��V,�g��t�H�6̌�<:�숄Uy7L��U���BSt�1�йp]�	UK���*P�5�
L���ws����;,i�+���T�ETm�#S���/:��^Vx��bT�0(��Y6��E�m v��ߌ����R�0����v/�[�\�*��C90�%ə�c"6��3/.Wɓ��v����ק+1�bGZ��=����D�����$J��!���w�;RKr
�#,8���֫��Tj���� ���+H3\E%2�fNXqÈ�9te����hn��/�puq�o�f��9�9��;O��l�2辿�j1E2%����h�:�E��vJg�Y�S����c꼇��ڑ,��J�H��y�3�s��ӗ_��LJ$�B������d<�z����Г9� #:!�����^k�"��O7�$G�݌��P��(ii�.}�]X��7X}␭��	�u���/e�ؗ�tfwI]��c���\���9���?�{�Em�� s/��D�mn	���,�M"M��D��ФC�����{���� X�@.#΀������0u��P��[��x���
a"�V=Lz�C�ܑ%W�zY��e��(��[��m?>���tƻ�>)g4G�b�{ң+�������!�C�Չ��koUx;/�~Ug�4��8�>y˨��q#��v׏g�b��&��7�������iD/�=7�� ֱ~�ʶ�Y�����N�vC���c{�"�$����(�H�M�HG�x�#sAf����p/�%6k^mh�`A�bTDA�S���3	��\�k��Va�`�:7�[6F�T+�,���B<�/ɘR�-����H�zꃃ�8n�U_;	��������⥘�V�y����f�0c޻m�F�u��xIa4�U��<A���,��h�� 5����j�]��l���:��U����#�_�����b̉^P�����)C�b�Ѯ�؀�+�Ngr��͋ ���#���w��V#�V
�c�D�mc+�sUk�^�RTb�@�G,q؋�ImC��zh�d���\����|�^9b������AѩR
Q��Y4��{JӸ�(Q�g�1$��@e�3Ceu<�7�U(��:�j�s���.k��/�ӊ*���ߋ�!��M���}���S24qÛl��#-�<���.�Ȓ��9��0��6�K}4K�0�K�����q>�lZ޳(�R��/��Њ�˻�]U_J�5#8����؂?m�������c��V2��).%�����pf���ddd�(�w�&.k��~�ʫm�������n�q���S(�{�ɋ�&*+�Z->�q��;��/�h���vzיȮG����j�}�{^����E��zʔrc�Z���;7G�f�WS�#���-A�`d�N�Ze��s?��4��:��d3PUd	
̟c�B������p�!��`Ԃ�"r�2g���Z|%��E:A� �$cg�
)���=�'�ȩkF0�AZ��������1I��W4h���N�e�Zލ�n��̀��2�F��+�4ڊ�`:$�V��f+
�僧�o�_F0~�:�b[�
����������C�0'Neή�{��jwX3뱧�|]4�w�����X�/��\��/c2m�nY<~�S$]��S=n�"EfS��q�v�~��Xc?$��� y�K�J���Q��Ll���)W����k?��A}��p�s���y�y�@(΍������fz�Y���VbM���&p�(Z�Y:�<e�'�!���ː�d+-��5�L�9� ��;�m������-;"�4�t�&��I� [J'�N�8���l����l�#F��mĖaM��Z��ZY]	���CkP��$i�^�6����\bι�qӤ<JH��d)��y��W��������F��5a6��&�O͙	[�b5K Z����g��z�^��������[Mxjgߥ�R�ks9.�e���ST�4��ka��/�m��X�2�A���l�9�g��;ɹ7f�J9�Z\��h��`�@
 '7,�0B�Eu�@[y`�}m��q�����a ����٥)S���Ƴ�"�����4o���}>��`�(A;[���Z`D��m�B.̀�)�;�w����R�,�!��RO�g��+܊eb+1FB�G��̋4c��w�GFe�r*N,%j�Rz� H*��m�Oڳ����e��v�V�*��6J0�h-F>�H�y��]��H�[�]�>A�r����C�v}\<���nF �g�1h�"Cn�dU8�T��3���)+|�@$�e+�Nk�ƛ&=0��`s钇JL�F
�MtMѰ*j`����G_�m���gE�)(����!��h��J���di������&/|"0#k�?��sz���{à4��c0̨M���פ�LÏ����aE_-u��ٿ��m���P{���X����c�@�ؓ@�Ȝ�q�bd�G����D���6ڟ�@�,�N��� �!�r|��S\�Y�:J�3���4^	�Ⅷ�o]:ֿNSm��Eo����t?�����CB%����n�d��K�n�[��A���4X(ׂ�lF���6�7J����G����� c�ل�{(��́�ȵ�X�/Q��J�3yO曲w�d��$1�����SF��f���{� P�����_�8Ճb�Gl"6�L�����pU(F?����l� ��)���wϷO�)�T)1�����kٕʦx�AnH��~��^�+�On�г�ܹ�/�b(���s7�CmQ0kx����\�a��vl�����p`��]7ɸ�i�c�b�,�����Ȉ�#�[{�7h'IQ(���}%��>�<^��R]�	&A���id���z��:mBs,b �r�X�|L���d�w�Ε_��20�R�6�� #������S�w��H�$��3'�V>8��3�LӔ�p,��Īy �������u&&���=j�M��D��8Ff�/����-n˩-�d8s* �e��gۇX���g= ޛ�a�iA���P��g���<�_��
T$J:2�,��oԱ{�EH�r�w,����G�GU�#L�1tyK(�`�!0�#�o�&Js�<盾�w��G�z5�
��K��;�5��D������ǫ�G�ل���VJL&x��X���Q!�@�O�O��Zy��՞��`�blw�f]� ������y�Q��ޱ[s?����C���'�ha�������n�x� ��]�A[W�z��bx��x���B$������nv�˫���q������W�3m�Q��7e��I�����8<��-�9������l�+D�%��}a�j�Ԏ���Nn;d��~�t��;*���ۍe��)����y�88@�L���H>�}�^wXb�@�Ǫ�����k ��fu�ȝɡ�e��4���z�Q��݂q����a����<ͣ�}�{C�4��*�X��Z�¿݃c�%T���jjձz#�c9���*�<��7��M3�dE��"��KFv����k�7:HR��o�0`u�L�j���y�s��8�gQ�};��פl*�_1�(��~r�
��4��������^�EN	�P S �����'��3(��\��'+��'ts��v��k0б)J��bIq�j>�(��CB�����u�A��F�i��g4���@�q��I�F��F፶�r��JlFV��*�=Vk����a�K�䑔�*Փ����ߖl]�'���Ĩ�/g��m
�]>E��=w�ln3Fi�p�_��?Qkz�CR �
���'�	<5��-G��
!�߂4�R;,�~���WZ!���/m��� JI�i_���R/C5U��$b˓�]�A�3 f_�z�������-�E	�+b�v��|Rx9%�E��[�cVdOƽF�KV\��c���?�	B����a����-�eJ�����:.��+�X����V����A��{���G��� l��0_(T/P�G�U^z3�,K��V�Ɉq��l��i���0s��b�K�8�%����g'�2� �%�|.Ly�1��RXX�?*���)�(�f�l��+����{hu8�e���l���3��֨K���(��Y뚬�xJbͦ,I�;#�J�5.���H�|��2Ù�'t7�$=I\'x*).�>7���1S��\=H`@�g��d�J�T����Rs�#ڵ�$uι�T�~x��)��	�+Ugqr}���	s�0um�-��$D�i�ǃ��^s����N�o�C�?��Vے�<\E�#���x��D����9�KeǪ�I*Dq��6�q^�l_Z%k��ma�����ƅ �[�0��:"��q��Ϻ,�=G���,�����l�ᶟ<o#y�J�W:HAt B���
��׺+yg�h��Ơ�C��R��t��C2�ȑ�ܹ�����eߢc���5�S�&�/	��^�Q<O�[�=2���|&��/�U��S�Ù7��5#����VG�}{x7;�}�y ۽h��lyh��	��;r	(\�˾>W���Cɦ_$l3l�d��I=B�P�J��)XL�?�%w�.٢��>������:JV`��t!Z7Y &�n#�c§!+�3�����3�~��uv����=��sq��&r �۹�T~�ſ�xj�u3B��+�gm�"�O������SC`���[�V��L��^�eA8��UC�o�\�,,�$�Y�����@N�/Å�AmA�I��ڶ'��������A�g�@�Z�X�3�L�p+��M�$.�NW�v^��w|.�څ6_�f}�|?�p(���H��cg��L3����;^4���'R:l`��I!�ي@����߃5�yo�����\���;�vVVzgd�E�t���k��8�j*�4���-�CnG��G1�r)�Nn%\!��4>�������$�Ő�tx�b�3�����i��p&���5�nu��}�I�Čn�h�6H�}�1�^� H0��\���b�x)_ e�����`����)��Z��ߘ���gP>&e�i"�.�DZF�s<�Z�!����v &������_q�x3��HF�D�<m�.��{u�~��ڰH�Y0+f�֢��t'�N���^[� ��]�*����ː 0MD��}�^B҇���b�E%W6��g;{j,�[�X��,̯�l�r�YDkQ�����ܶj��=QY�3��9B9��yn4�F9{g^
��@��
��k��ң �������I�<��DcGY��ʚ@#����\aeDT�8h�����Ԛ<uT���z!/��la.��	�$�e|�؝��#Mh�9���l��}q�o��#a��l���p�E+��G%o����t��]T�@� �c�M,n��N���s��2n�-��T�Ko����v-�R�B�媼��{����QÀ��	+Lht������6�S�}� �S�L�&��5a7��;%�hc��9���u�^j�c%^�TnC
�aW^�Rh
ʶ�k����KQ�?e:a��������;nT�	vj�(��f0FJ�h���x� Ɯ���*�r�oF��`�S)����7"����/�ޭ��0U�g@�Xa��t�4���1>`cq��񮺖�̛͔x�_2�\���	ZރW����tH�=�� ������`�B+{`���)]sj�X�Ϫ+W/��w�bP��@���#�Q�O�2��`]��K/��}��O/&SNx7˱L̻�1�L^խ��t��(;�V1�̱�:�oO�yQ����t�H���0h��gutk�D.��"��-4c�ˡ�qg�\K)ls���a$>n�cQ(�޷.��= ��R��cӗ/w�z"�`�����ǃ����dW�ꯞ���	��vƢ�S��nCh}�x&�C���zÄ1;H�1�i2hRY6P�Ω<� i��Q���D�����0̼�M��S��e��y~.��N�[W��3��L/n�!l������3��o�K�s-��4�E��{#��X�ɤc?͞]���he~;C"^"Wd!���%tO�lZ!����&������uO�@�6�sj�o�SO�7V\~ل���������l[
3��隤�j� ��4��js�
�ℒ�shH�'X��=�#�ݏ;9	)0�赿gr�u�.������ʍ����d[
�j��ܼ���&���Ph�씜�	�>~���D�{~����"5�$R��B�}���v�����x��
��Û4+R��i��|�@'��ȫ4�H�X�I��8��WV59��gl��pNdq#n��G��	 �'�ˎ[�:��G��֠�<��K���վ���Dt�m-|�He܍���*�� ��ض��8Y�v��\u�W�U����9є��Έ��kf��sPv���B���Vmv����ܬ�p��`�b��R"I�"��D�M�m|�Q4��~��BH�ϒ���8?k��l8��~�#�,���^�8�j���(���xZi�� ��c�q���e�I嘳8������Dl�V�ZF�e��b �G̅�Qֹ��!1��;�8�!�?����7�qo�6�~�	9�}����,H���ǲ.T�Ϗ�Z��"�/jSO`�T�
q��w��y"�p�k��>�I�=U�d"����_b3�)6�'{��4(4�̊�\u�������&�l����e���P�Į;Y�/��s���t��<�v(+S���e����ð��F��n�0�t�bc.
�jY��*���CĘ�Y�骹��;��م`k��!�[�>Q|/�p��^���S#,,�#��x��Z���@Gc�GI�����Q���e�ǂȟ���!�J���$�)�j0a�����^����b�Ώ2�Mt��1�#��ÄR�����&Ь�q���l�$'�o�J'���U%���G=]�ܧ~%�����t�8�����E����3�k�};C�Ĭ.��I�ϫ�̦����t�fm�$t�垌Y�E�A��,ݧ�QH��1�_�����v�Y;��� r�L�)������J���跴a~�Vn�j?�j}#���}��am����\�������8}#tCH��:%�}�@q���F��^#������1]t?����1�x����2��)0̼��׵�*,x��W,0m>��ы����[q���)96��~�T��[f7:����i M/Q���۸s��	�K	������t)����51�%�iW����L}���t n�,��~�b:�ZF�7����#���,m�������l������ ō�$K�G������Z��=ߏ�m{L��t�5<����o������@w"Ri4ߍ��3��A���TY��L������0"H}��OɆ���1h�O�[��v���|��ָs,ʅsx�V33	�&̵�웲�c�b5�U�Q�9���W�9w��۽J�h������dB����<!ǿ�\*n��ia�k7W���qڊ{JWK����c��g5̦A�},$�����C���Th�V�qQ Hh/>������ъ���"�o�������:�`Q!y5��K�`�N!Bs'�%����F���H���s�Ջ�L[9�]㶱5�2P�O �2���ڰ'�>����g9E�-R�!���/�� �9	��$���w��i���~}9�b��f^��ִR][��{+CB��[��]i֒�O��t�k������2b��Q͕�?���k��S�9[��ϧ�~g��dU@�z�<l���)�"na�r�=�E���%0u�����6{{w*PaL��{V���|]ĵ�g��˭��@�pz���8`Ͽ��?|����I>h6�<��YJ,�u�d�\�`տ����P�֔""܇x�&����z��B�pj�<#��Z�F���E@��~~suD���s������/𭖯�!�Yz�[+l�#�o]���Cx�{��V}G	�Jd�&6���:�W�]��"jz�����6�3�� ����z�x���+����������,8[_�DR�6N;��I���w9$��8�|6��6:�i8�}�nYK�_w�o�%�5VR�r1�q ��Q��4uQ��`c,`�o�ЬG�ޜ�m��Ń���G�gNئ���d왨���9�X�X�`U�v�5�cZG��_-��]�n������_S7B�*�8�f�o�Kd�3g70̾��k3u���Vi2������'_W7��e�8L�g�;˙�q��Ȍ-�X_�m��׊�KJ��s�Dñ�q����-�����N�w��ЀD���J$wy1�V)2	�g���Q=iF����g�d�B�&�>׻�d�/�A!�4��B����2\dB���
�Dn}U��W'סm�Ԩ�!�yt7�`Uy?"|VQ�ȡ�p�k��ꕙQB�v�fN{�L��NGqڹ�j�p�(�͏.G��?���c��R������c�X1qQ�ǨŻ���9�K�yyN��V
��j���֫k� j��F���C�9���X�2Ha�Pf�L�wuzj�Zr���7���T��Xg��d��
�ce��-w�e�_S'��V������[/��*r����ꈂ�����̫ &�!
�V��^�@�j�$n����s�}�`_Ү-�?���v@6$EVe ��3���H�������Ř��Z}�|��|ퟐ2TH�:T�V�Z�i�.>�)U�q�wp_�2R���=f��Y�ӵs']Dj�3t֛W~�[#�t�ɖ!,�`*E?�`��G\#����O�{�N��'�̀.	��G���ӈ�?�fR2U�]M�^2���ÂK$?�ت����}پ�e�ٗ�Y���]n�,B4����{�&�^�U��
�w�&D7�=�6��7:���ʒ{Jb�H��6�5�w��>�>���@�n~r8�Ps����:]�N�)<P��*�̊ˮ��`s'�,k!Ԏ0�桾�Ӧ��I>:��z�7�7�N9��%E5��X����$�j�i�b�7�{��NCl�x������������.qC	��_�/A2������+JВ����rK�u.�SP��n�3q}ۍ-�U|�D�ob(�磍%�r�I�ܻ�O|���{�k�)��d7}Ǯ�/}��O�k̽���^mg9��~���xV��AJ���N	�6 [Ç���0��yH��U�^�1�1��N�,ޕQ?�j����7/-v(x�.�!��mA��(�C��z��O|@�@�ׇ���@P�rD}㰏Tv��<�o�2��Q��>D�"��c�Q^E�"��Ьr7P�i{@�F�T�R;i�B=�Ʀ��
[��n���%��uV��P7Ĩ��;�lC���xz�\�C���lxߑ0���h �hd�-�D��pl�ge�fQ����e���`�u=��	�kVϹ���i�G��*��>x���VZ��2B�ƨ�d��f-�*T��|	��A)g����K7��x'����#Mv�vu��l��Җ��dߒ��jǇ���ܚ,���o����a�Nԅ�M�1Oϯ�=�:��9Aj7�fh�$�������I݄?j��9�Xyb�^�'����V�JGj	�H�־˅%����K�3�F�꧉h�_?�S�&��y�����~yNGZ<��e��M",t��f�޻�Q�!�В�đ,�6�;t����$�=z5C�����n�˨��:|��h|�.~������f�'d#/~�4�Q�ad�h�ဌ��*$g�.����m$��`���H:��	�|�+6_�
;n�\�3 g�7/|m%�s蔅�69"V���}ȞȽj�w%��8�>Ku2��E�ԏ��I�3�O�Χ�o�K�Q�r9)x�:>�� 8����Bn�f����g�?L�8�:'Tx�����3�{��⁹<CǊ�J����G*8�G��y�Q~l_�c�Zovx��H\��u����i>���u}$D^'����sT�^������s��֏�aw^(?ށ���Aԣ�*ش%�[w&���E�Ċ��!m*�#�x�, j�P��b�0Ǌ����̝k��;t0��J�L��X��pY6ǫr;bn^2p�&�F$����ɴ�y�R�	6z��1�5}[3;����xO���D�p	�hO0O%�2�ݫ���dK���^�8���8���k������cl���)QD���գ����(�W��z�m! �{h��zS��n쁔�{�٘�Sl�5���k��: ���R��F���YbX�c�a!|�.K�d�x�t�:�͇?�U��)	gH��#VǜW{hN��t�F�����E�z;�B�c����TxU�� �0�O�d�\!���GY��d���ӽT�;˯E��g�{��Z���=��-э�g�9���a����~fᔛ��hD����!+�f0o�9�A~
NPY��j9��Oj��>�o[�8�a��"��l��[�L�z��Ӓ]�Y٤m$�B��]�[�X�Z����Bܞ�
�æg�H�asg�5L<�E~(lX�y���6럏,�duh�5і�#0��H_�j��G��+"ׄ�Ӥ�i���}�j��=1�Q������p�����atf�k�ni�0�@��F�v1ŐvdɒR�@fy*p~�����XJ���{T5��@��j����� ]+��a�&��.��Yo�������ӡx �8�x���x����wO�*Rs��_�w���	4�̕�o���e����g��Weھ�L9|�=x{���,�vА������ǌy����-�JU~���N}K�w!����v��SUΫ�)|iU�ş�f��	8F^A�uኁ���FL���9U��h��f���1��
^r�)O�P
ֆ���Q
��Xu;�P?|U�]Z)�%{��(�AsXJ��йv� (��z�H$�s8`�Kqj�k��f��6�?J�~ڣ���fp�&Zv���/ ��Z��2_@a���*;�D[�b7�Ƚ��|�hӔw1�6�`�`=�0�΀�#�Q�G�=8�{E�lK��Ө�OK�+��o�~Z�����6�������o��]E;�3�]z�8Q��N L~T���U��O����s=�C�x>#�D�p��"(�>�Z0�D�I�k��*�x�%��ɛ=���S*�Ky�Ǣ\b"脬�7t�.�m�Z�	��>�:M�t����.��L�Sx�pd��L^Ȏ���H&Dz��0`�5('���+����Ɗ�-/EV `����˕#����v�>��cD	hYJD/��#�����'1����i�O���v��$�s�Q�O��oE�`j߽���;t����
��o�;�푖b!��`b��>�+�v0��_I��A�]],�������Ԧ8�=4zMؐz�X���hA�o!�E��U�j���h��V$C/�p���-��B��g�W���,[�>�3`�2�3X�
ǡG#�q-Z�*�7���7�|�S���J;(j�L�o���w��7�`g�a��Eh
]����̭�ۤ	uc>p��(Zk�ۦ�Z`��G����l�t%�maө�DJȀ\�y�TSD�E�i�搗�H�1��VX?��W�U�M̋e��r�ms��$ߍ���_�����zAWjJhűXw��o���b(�H(8B�৳B�I+;q���~�+yv�?q:���y�¯�u�d/gz�&���"���� 3�H3q 4�a���6��+���7�����$�����Dlv{}�L�C���$)�e�~\T�x[��=B钄�����o�wbS#A�G/i����̺L��SL�߀{|V}�.u��L5��;�ޞ�R�JH/��&�WR�Rk�4�
�G�������|�H�2d]�c���g:~�C)�>
-_a=��3��e��=j�2���h���￴ڵ;ʌ �����Nj_^$�2�/I��9F�v'��U��ƾ}Je ���rĢ���%�%�x�j6��i�� #��M����I"�l�3�P�9�ޮ�Zxb�����?ʢjZ�͹^�Ur
����(Q�L ��5���^�����H���"m-�N�)�l?Rk��m{FHoS"��=�M�����pv9���SJ!��E>�p3N�W�ui���('�qv�ɰd�����u�`�t��8��Z�ѢT�b�����).���Ŧ��W����3w�O���j�Ve0�b��q˧���,�C�rr��:2����K�~P�Ԇ#�
�D��pb-SŶz�iY���l��JeĻ��Wp�Rl��=h`�����`���G8�ў�:�4v�b��p�@�a٣�}�
J s�r��9
I��x�����f%�D�9�L@�4_Y�֥z�^�V��o|nF�'�ً���8������b�'�1�UJZ�L���|WM���6�DX[. tmy�[Ɯ|Av��D��G��S\����p#,���iǸ����G2��������Qmd	a��tH����ϜF��S��)���.t���X�qG�T���.�/D����p���s6�߀�8r�������Ϙ��xȼ�e�������.�$x6&�P3�����m�Op���jg����y�l��c\��ێ��!c��pۦ�5t�_�E��+�͕�ǗE�g�����Ӕ-�>k(q�؀vg��pS��2w-Gy<�X�s��X9&	�pq�H��`�[�T�	�7	��I;<��+��W��� �q��Y�����/�w�U�H)P���\>:��Mqw�Fv��X��Ԃlt˵�H��18�V(g1�^!H@�ŷ߳�3U�(�8��J�uzs�1�-�'�Z�if�F���4l����	�����mq���[���K,J�U��qڥ���y�г�����m�w=e۞���*��EV�,����jz[j���'X�������݀�"����Y`�8��Uy�e��T_�կ��[���Eʰ��r@��b�5�^�gAv�h���Sn���<��r��6�T��#F�������f�sW_a�|���ҕ�~8�%e�C=� 9Y���sb�S�M0����o>��d��:�����uQ3��n%������'HT��B�^���`c�=�(�S*�6��d�Y�iã� u;�^�J�@��0�W��L�n�W�AZZ�����krj�5��<m#�s׬e�lg��Zs���&��r|JZ���.n+��[��?%l?���`E*�"/P�G�Y�0e6v_����K�x�����b�OT*_��U�����]�U��ߺ�Vi�*36��Fl �4�j�]�q�1[��M�Q���K���Y	�%s�3
�F`ೳ7BbԳ7Bp����ה>�������֗�n�4�"d�ɠ�Fe�}���T��t%��aT��I�u�#=a��TLӟ�'��&��~l�d�s�����j������]:���҄�(ǐH�Tn�̖1�_�HWզ����Z%��1P�hD��׶�T�\�hA�,}���;}��v�L�\Eݧ�m�O����ъ�><*(I3l�|�we)/M� :֔ah�(Ψ�Ul;,Y9´K�H�<�m���j�7�ھFsofA`��~Q¢��n�-���q�(C� F�f��m,m��T�
��Q2�~O"<&��ۺy�͸g*��s�|(%�ڹ��鎍��˿?��fəD��?FqB�	YY��a�jBb���S~�
@I~���"_����{�h�����h�n��Dx�$��\#%�0�q����������W]L�����=�����9��>����?2rɩROf����I�l�d��)��hU\�px��*B�uَo֐�w����)�AE�iE	������N--XJ!z]J�:��}�(��g�aA�r��U�xb��q�B��U����umWT|vh�Ɉ��ވP��Z�!<<f~"Ot��e��� P�� ���e�U'Z�wĦ�/m�[�Ff���=?�n�j��:×�������ಠq�9��No�;u���N���b�q~���ij�\�!�Cq���������=c�T>1���<������kKX���@����F�>�IQI~����\�6��Ť!$�Wɲ�`�`��B��gx���i�W2���uV�Ƨ���{�����8�#�LD��LٻJ�?)V��n(���c+�I�����}p��1p�� �c,����d�j"1'�N]l�n�H�oJ�g�ƽ����|D+�V:?V�
q��u1��?=3��93o�(���p��Պ�_U��S��D[��Q��jì�/$�ț��s�g*�#�XDu����,s���- ��5�+��q�1/�?N�gdqS�������TK��i�6��+��05?��@���G�X����sEg�v��X�Z+�0GbN��&W�79GX�uKŷi\����dr2YtF�c�X��<�{u���eu��D4�C�ev���e&�ƅw�_��~�)[�C)�$�n�p[�* ���@k� �#-���Y��vX�����N�
��LO�n�H�*dUs�*��"��'䣺cc�(T8�&��D9���j����7��?'�+z�`-��'�o)��Q΂ӏ��y�}nRT�b:�|L�.99�ؾ$;�U#Ú�}���6nmI1�Qa��P�fS(�.���1B9�a�芦pV��	�GFgjNN�T�&�)�kt��O�M氵�թ l.#a�eld����]��L����I���z��Mx�K�Vm`uQ��+6�>�(�k�˄� M�B��^�w���8z- D��ru<������Q �!����5~N����fw}�"!�o��E;f!�X�~0��j�<����������$#�hK�ĸ���0S��f�*�F<������]kS�wLe�&!�xRƭ}x�ԯa����t�s�Th�����Rۋ�ğtHH1�a=lrL��sM���-� �GA��<�y���K^���b�@����e�>�
��&g���̜�_�z�A$�*�_o1T�<���x����2��y�xʞ�%�[e�/���pC
���x��%�ujk�*v���&W_Z?���x�
�Hÿ��a�� xZ��)���btO>�����,���1�ܧ�ĵ3�i[��t��{�f�d�^��3@l��Χ��&Iv�S�l}�����3q��Ht�r��Q���
�ř�0ݒb��ݭһW]��71����N��{��XJ6 `.�b�d.н�!g��%z��H݇�E�|Q��(׼k��t���B�k8�e���]�VJ�F��
����b��8?ܔ��*�u�7�#X!�m�x�q?WEҿٜ�y<	�q�c���b�ʖ�Crً�:���}��С�pg�d��#�=�=/��(���s�7/:\Z���@;m{��p���Hs>ӪtR6��v�M����&;3(X�k"d�JtA�EZ.{���Y)�7!�^"D��bp�n�S�a��8�٨a�,@zC�f�ø�=�B$�b�I�mP����&�+V�P���f4}����:��{2_���,'^#|�n!u���8+��\�Vϛ�3����{�]��K���S�\��A:�����=�!H&*6�m�;�3��Q쒜ߦ�j?���&zp��s�{��-�B�l'/u�yǫ{�$���4�Ȥ�(�ߠ�����'ח��$b���/�f��{��z
q�����֢�3���}^��0��g#Jɴ
��iZ�@>�:�M!�I�����z�����,#��Y��N�!7֦	���6�F���.�CH��*�����1��\	"��W{��FCDb�pz�2���B���Ͻ%HI
����*
�I��OS�4��WcnD�1�c�m�+�N��ċ��z��H$�}jv�k�u�
cB��V�/�	g��1���6a1��~�Q��`�~=bK<��i����V�:�묪�P�G�o?J\�Y X_��3ڵ��[����X�Ӡ�����/z%�Yp:��&� �����Q��붏�-�� ��tź��ۇK�^���>�(��˒5��#��D��a2���^µ��4�Ek�f$�PM���a[ȼ�G�Ї����r)�0�B
�)H<�����_����H#Ix��c}Q,��צ	P�3=��!|�O:�A�/6=��H�X}�A�G`�6�K�{�C��W,�,�78|�z�������`I/[>��������)笤U�`iBJ��/�״j'����4��������#^W�u}��,m���C���յ�8U3�kS� OYm�|�v����G�n0�~ܿJ��v����s~��ݔC�@��J�]K�Qvc�S9סA�ܵ�V�����^�Ф�	��6�A�'��1��Pzm`�Y=�fH�+F��L�[��2U��	�ZJ9�T��j �޺��������ڣ�����>)�s.s��r�T)��[�b�K|{���|�+i��=��5�BC��R�_d�9�x�״��=��#�N`�ʝP:O�T-nɼ%����lǣ��	0�h�.}�
���kA{�\6���]�4hRAx����6��| �,��|��d}U"�~�D�gć�䒴��M�uZ��;u:|��F����55I�f.HZ��^��Kb�A�j*�;!&+NK�L�BK�c�V/&Ҏ�W�n�wz�T�*ٟ��E���YA�H�6ǋ*V�XO^.�SM��O��3k���ڈ<�Uzf�d��
#�g��`��,��%�{W�Z@����p:dP*B-��4�I�D_nu/��̗���N0��^��_N�c������ύ�K�12L_}�5�+����u<x�2x\{<P�]2�w*�xW��ǁ6@X<�y��d��J���^�!�=G�]�|&ٸ�RXm��]���Q������.���`,��7�E�`8�"�kz�����1e�Z�!�������7c�
�
���85���9���N�o,j�W����4��ب�TI�lN�?M��!���o�f�i��vQ�K�����Ė�R�����L��oޓ΢�l��8̷`�����lT�
��0�^(��JM�)�xv+Γ�h����q󮝂���2k���J���Rr����bq8��Q-8��y� ��2<;���O�,7�����4!�Z�T�����R�ڒ�ouШ���3T䎭�'�uD�2�Z�=���n;�MƩ��n(ˢ���2S{�=�0�c�w���0C���<�v0��]�2ˑ���Ve+`y �4,�w�T�Cr#�]�����LN���_�F*���[j�⹹*���T�V�KF�l��R��ޖ�U����h(���,�P'�b3�E�����oߊ��C�6�O]sBÁ�/m����_�5��q��֮,�(T�S:#����z�.��;��y�J؝JC����z#B��rh��mͳ�1�ziִ�EN���L�)(�L
�Z_.�89��?a�7�F���A!�-��sa�d	ma�(�q�4��^��?V��x����N_�?Y��y#���Czt�V�D&�n+�� ��=���t@�(���N���#x��!g����W7l#~���O%s�P>lAW�*�����L����9��y��  6�.h���ӛ}f�V������Re�ߖ����=�w��j�/�$���/�b�����I�	�G(����eo�O ���<��J9�y7�ϓ32xN�$m��_u����P��H v���K���ns�^գ�%�$2�h��Ly�)'!��}�]�G=q&�Ӓ	�d*V�K�P��9��$�(h*0U�vg��r���:�ėNwUzc�Wl�.嫿<}�U���-�Z�J	A����M�����O� k`D��s� 1�h9�Z�c\}`m�T������&����!��ى�Gm��Z�&�`��&�L�M9���� cQa�:!T/M�,'����X�	g� ���V������( �\B\��p4�����v���Vs>���m�11�ˍ-�s�X��4HIӌ.��ի+g"�Y�u�)��ި4�s*�'��9��rw��S�֥�F����.��+?�žԶ�X�{]s�<���2Qh�_�Ru1�Wq>v���P�R�Tc_��CM\<�����)�� ~���W���͵���篞,	^��@v���6�ބkƝ���-d�,`�QV�U�`��v����֚��[�nR�>0-6�M�l}=�)�R�ѽ0ŭ�����VWF��`TS�kM�9�����G��Ŏ���;����B2ۇ�aHgZ\���,���g�͉4$�QwB�G�'�*y�ō*��qLs��"MW_��~�X�{�f����X�rg4�)�c���8s=�]c�l4w6.�MP�3�c\]�y�鄗	�hG ��R��zeB���p7R��	i�-�e��w���� �|�� ��$�Z+��p]#14)~���~�y�q�wA,�����S�d�Y��-�_)��J��҉<8�Z�+q�۟�5�#�kG��O���|��~���3RB͘�����L�kg�q�g��U#�Yv��Dv�'i���.���L~���:��0�:�i��"���W���|���[�WeZ�I�
��_<2�\V�3������F³�-Qy8<g�2�UdK���Բ्�����Zי��.��!|���+x���v����K2�%Bp�=�SLßG�������S<��� �x';d�"i�t���u$�i��E��B��u�߶�+�+�׬�D4�Ct\!�7�Ǥ	k��z/q}�Ț2��"�#��<޷E��
V*U���%�Lf���.�@d[��+���7F+&kQ�2-���
w
CM���6L쯨̹4��*�˪�Ѝ��p��0����
���4k5��#�]�w��'d�qu����+F�a�R,���&A�̗�.$�/[+��t�'b�:2�xRݷ	?Ӝ5>�<�PS"#b�C�ql�(B�4D�Z���@��(V��׶�HBh_S�{�xL�B�O�¤�<�x�d'DQ�5A����꽹���9^�� =��w�XJ�B	c1~���>n�e��R�b&��P����Mmk��X]��wq|�j螼ڃH����ى��h�܋�:����8/f�����uR틋�њp��}.n�:lI�����Ƚ0^T����b�ui��l�& �I��K�9Le+���ٯ��F������w���aז�������� O�� qeK�mY~8-΋������ ���?�]�:P���7惍J}���y�"@�Y�(yQ���r?跜��ϼ͵6�)�U��3
=YW�w!����t��>��u�����2��Ҥ�Hj�K.��_0n���$��K �{�=��(�͌V~.Wg|���P=v��)n��d0f��g��\$WP1��P3��"��Y��Rͪ[A'o|5�h��0���`�j=� L1*z+�����|N)��d7��]A�=؞��u&��m-8:�M�J��>��i�8��b�|��>4R���S��|�v��̯���[�g�mq�1O?�r[5X��σ�$߿{�;��q+[[p�fk[Ӱ��W�p�y�%[*1�VUGX�J��>Fk׮S��ioM&�E	9c^��r�B���FF�΋Z'��D�'5�d;;������X��t���rp)o��2���#_�����E{RD���"c�����f�ʫ294^��v?��~c�@6���7�ǽ�Z��\QԹI���wV�~n����q8h`�H)�����&�:&
�IT0:����|��?����(���B7�
��;?�޷�O�Nn����?O������Ifs�[i`s|��T%�t)o��ӏ(���:,���cq�<�rx~�ҧ0[rǅ�p~)��^�XpeQ��?�'����,�U�rPp��|s��@tE�	Ԝ��������I���DKkC6c �Q t�C��:VCg���A�^{�q ث���XL�����mk����bY�wa�e�ȝN���K��)k�#2V>�,�p��Д�>�-5�D���6:o�uކ��#G�������1X�ͭ���K7Ъ`8w#��]U�K$��cԎz��"&gatkƠ�${�=q�y���75��#����u�h��[��?s̢��G,'j��y��~~�[�T	>Q��M8n�sK�h�F�6Y��L#�2�E�:쀗��W�"���b}�u�n'S2N�F���{E�v�gGDVy�n8{�?��o����~E���y>�a&��0Y{��S����2 [���IU�=6�W��bH�{�(;b��K��?�>��I��5�|�Yb��ZE_,��X�,��w�G�M
��)ݰ����n_��It� �r˵�����ݞ��y��+��F;����'�HmB�R��ҏ�%�w|�@�a]�A�Ƣ���<�H
Swp|��4T4�`r��8f��e��<���E�&"�NaRƅ���:�!�С�j��X~�ߓ[�f���Fȧ���X�e��6Y��F}��C�u4�QSZ���Xq�Y�ӓ����2*�;�t�b�OoYp/�nFv�����%Za^x���5�SO;�Y�JF�r�~�&����6Um|��^����A��8$�GMt��ΧNC/�+l��3R���X(�����C�<2L޵Y�D;F	X/mR�;�c��S/�����Gg=���K�	挰�.�|\����AP�@B�ɏ�bO�||��K�_������ȡZ#���ц����C��`k���:�	H�<���f-Gn��#�ܸ5�2��#���ބ�C��IÕ�<]��Gmx^�K�oP�M�2�l���������܃-b�" O�U:y��m��}]��B��?dVU���y�̩Y��x)���=�A���V� ʙ������v�l���:�\DΤI�!�����9P,N�`�������A�z�]E�����N���֬��l09YJv��L�י#>�/� �f�Q�R�5�P�R��{��S�.�>5�T�d�H�8�_܏�ȣ'Z��"��y��Ŀ�*�q:�;n�d=`+�	B����w˻�:��j0D��:'O�].�j�"��CYQb��5D�y�2[�J��e����ӻ[��.	_o���J��̺�kl�p�a��k����ٿ+���r�[��5q3�Z�U���OiY}D)�������Z1�F���P�w�ڋ�{�N���"x7/�M)���7�m�?�И��Bp:�K�D��G�8'SkBA��,XAI��6-{�6�Un"2/�b��%C4�n�~o�.Ł�X�6a�1��F�0#���-���	K�:`�A��!�*���������7iL��}\��dx\o�O��(X�O�/�6��Y��$�F�V0|�O����2`K
8��}����7J}�����j�����@֫BK�t=�i�����/��������
��n�Z"7}��N!�d�9Q�׺�
��-�D>��c=B��s�՚-��Q�tSU��ny�������^���[9�����-��G%bt��߁kV�`�޸�u20$x5'����s� �Z�D�o�͎��䱩�������ϤY���`;�'�#�T��wf���HԈRݞ�,%�˓ȊHd�T s�pf;��#5U0	QN��N� �ϓWy��.�v����<{w�y�E�޿�'�.���煆)p�t6���o�C��,��~ܿ��0��*� ����5��G��̤� #xkH�����-�ɪ7��XHuPmt�Z�=�2BU9��Z�P ��ҜK��N[5��+�C��~j<�;jt����9g�f>����Q�����z� `L,z��Q��(>W�.09-j�q�t��5���&��1�Y��eK�`����Ӯ�}�_گYLT,�ԉ_��%yj8�X�\�Ӛ�I`6����T&�댾�"���9��2�.� �������A��~�'P��ɓg�[��-�Q��� p��=�����W�mP�xKG �8L�����	���
��u'3h�I��D�y	�2���]4]e�������/ѻ�m�&d�\��'���Z�>+c��`���9:�?!4���xƤ;�R� eNW�����M��2?�~鵁*�@D��r�� ��!H*�;��a��5��@j�.B�3HB�tal6)��o3L�tכ��m�����?as�f�?��2�dd�y�/��*ߒ�v�`���
�\�r�K��%��I���x�m����7W�ͩ.�}`��k����"Α���Gz�5�����RWO-���=hz<���`��R���4�]oG1�EV�-QA�!���@'�����M8��Ϫ(/��J)I�i�[��/ߏT�`K�"�E ��O ��"��b^�9RY��%9R��om��Q�9��ʹoH��1�O`,Ƨ�%v�]\ ��՚�y��ܜߋQ�M2�7A��H�����n�g�̞�ќ�i�|�0�wY�y	����L��9@��o��+[����˟5ؠr��l���|���z�*�'!��|���mG�$�Z|�����C�$�����'Ʋ�}K�ْ�/��Ia��)/��@B'JDq���~;��.�.����f��NRw��_����ŵÍ�q�\t,��y��� �Z/y�r)��u���9�v����_	�].D}�8�N�6KT_ݻT���}b��MG=�T�	x	�����=�j�g4W�+H޺�D����A��4����y�X>1{pNl��SI�`���6L9�߂�W��wF�ƻ�H�5��{.�\��7!=m`��z����'ԣ.X�ڎ��D�Й���fv�,�k>g��s{��}�c�v�R%�y܏>H��_̉P�4��p��\Ea��#I�o#D0�0��#���a4��,N�+	�
`�6y�N�*Z�� �ɽ�;�����&�x��0e���Txb���A�fQ4dn^��
����8�}bOn5��vE��چ\��Uhq�m$�3�Mv��5��&�O!@��*E�- �
+? k�&W�k�PD��݈>�����o��<�Mso�#r���E�������ܧ����s�қ.>hFt�>Ԏ��.��1	wO��w���,�B�Ά�dk�m��f��.�z�q��
�I�^ǯ�J��#$]4^��A�����(�K�Bj�||^-NX�(r�X��갸(Ɵ0�Ģ�Z1�}���>牖y��±�U?�Y�XDxF�h�8c��r��o��;�b�͠Fľ��iVF'�>�fU��d�$}$�}(�4���8�3Z�%��X�e¤�� :��a&�W�*����Ш�u��͘
i7�J��)9�f(
�'C�5��=>Mr��<��*ξa|����"�y�|7ތ&}��V �����O+�s����4���~��J$�Vr�2�����"x�Ɓ�L7 ��h�P�	A���sQ~�?�W� ����W�=1QKg�t�n�蛎�s[ߓ��.���4�)S�L;���8\ۀ!�?�|��(J�r�׹���[��{�� ��.��2�[�.QI���^mR����*D��U!�˘VC&_��P�.Y<�Bդ�#1��T����=��+�fYp8�!"+�ݤ2����D6�{n�1#��)i(U��Q�6.%�_�ߏ�Kgc���+�,f�.��
3��l$㣎x�&�A�"u��΋�|_��-R�ٱ����O�h�+w����ԓ��i������Ih��A�u��"H�(v�:$��tF
˙��+���,�:��F% ��p�fhȼ&��W�@,�37{r�of��.���$Z�M���6�*�l�[�b�)����U�b���EF�[<�u��#s��<��<*�|#g.�㈆�������%۪��St��Y3YAFՑ��i�٫jدG�m���fAVJ��)b�)cW$c�� h�-=��ü4�w���J�Y��݈I����omS&C�HAoQ:]-u���A^����L9����_ ����iS�>ہ�U��긠��(�pd��4��"N��۳�ij�~vi�1�?4#�
�. ���L\GbGMh�U�X,w@��>���Ȭ@C����D'�tw]���$�S�
��~b�ˊi����* ��'�̅P�\����2�V9�aE,X;�.�Ό]�����>�����r�� �4`��5d�$`}y�BEe�� ��XT�M�R��~B^��\Wi\D��_��-��M]����1@lq����-�]s�ω���7[x}2-_=~�̖�9�0K�1V��̸�ąBE����!�9.W��zC\��}�g��B&�ڡ�qL����iN�v (�M�l��mM�0Rs���,�X	����세Hd٬�g�G�Ir%T�K�}ë��L(�<�� �.Qw+V��d��h�V��oK�����f�~��g�ԼW��/���5�lN�P�8��	�ִs�"zD	8wńL�;_! g�M
��� ��.s��nӏF�A�{
I,����W]�����GkcȾ[�wuoaX���Â�2$�f�8h�~N}�cݽ���/��E�f��`�
���QR���I&iq�@zu�sr��	U�kݟ��$!�`-����nVx�)�7{�HQc�.�����O�p`�e �@��1<�KS
\��@�o�0;|w���}��=�������: �d�,�@]��{{&��=^T��}i�;���QHY7��M��k0qFg�7��7p_6���`K]�&�L�H$	��w�#Md�sC��)7*a��!x^�l�����0�������x��bJ>G��gȉ�ᮒ0����,	оEL��"��U}���5SS�9H ��j�����w�� O�vh�x~\���:]~&��O�0���v�������ҥCF�_�j�����8�,�h-Dz�|	�H<�#}إ����ش�ك@��0�*)�<�t0Y�O�(����1�8��G�$��=���� ɒ	����В���L~�29��U3K��I8Zڛ�.Lw:#q^��C�F��FN�i���et	�8H��_V~ݔu^N{{C��%�e�Fݠ��9G��lW*�s)����8�b�(��`���x��*Rd;��z%1�r�\J��^��BF}�(B/�x�c3����ܻi �`v-
/�6ŝ������nx��E�nE�c�k�r�jw�j�뤐��
�x��}Qu���n���Es�)ǌ�C�����(���l�E26���p��e*��[敺��u9c�N��M�q���/*Z�O���L#Xi�8p^n���w��>�����e������!�1`Qō
���8%緹�#��HX������-��(�o�i�#��C�? f�)ex��,�d�~	"ⵢJk(�75�˫2f��c~�01��P����]�Y�Ǟ�w�z�(T4����^'��r�g���t𛇏�́m,��7�����4�<o��J:I&Yi��/d%wG����8�w��Aեm_���fFk{`t^dHJ%�r�h�R����O,�t��M����0���$�uv��%�8Ɣ*BrJm�_'sml������Z��R<dǮ�UJ9�y�z؟
�yh�8�׀�t����(ٻ��g�МW�������?�zV�.����#�*��WE�lO�ԂʥM����p����l��W�0�:�o�?be�vj����*�J�O�>��0�8��ޠ�j^���A�"�f'��l�Ⱦ+�*!vK���N�^�9�Wg]��2��<�*_awjk�vq#r�y�ױ�̨�#�&�m�s��S�d'�h��	h��^�ͤ8�~A���&�F�+Ҵ�J��&��M�4�Y?�3��p���1�P��Do�z!��{~�U�K/���� ι�NeN�%��zNh�B\����gݗ�GX��+�rBR8�F �O����_���z��;�+�|gS��"��z�I���ۍ{6Q��r�:
�)[0P��U]S�33Z���'���F)+j=Q&	�ܫ���G���
��~ٻ˝А\�8D��U+�2"N�T�W��ù\��Aw��u-	We�^ѡj��ԙ�G9"Q�Z{:��S�m�>��jM�@�<~��K5���j		zbenԛ
߭I�=����eۺ)��L�!.�X�vb3����Н ����)���`C�76�:-#%$'��$����fK��� ^�	��t�f�Q���>Z����\���I���)�,e�Q�� �����K����G燓:�`��j6���O)�vP�`Qޣ���X�B泸M ��v��WY9�������Y����R�(-�O~tj���}U	���Bic���o���,m�ƨ�g �:���sHJ�n�&D@�?�er!$�Uz�!:������ǳ��X{E8t��*�O)�`�8NȦ
ĻwQ@��XR%��1C9�U��)5ohC�m��l������-nB�,C�j"ܑ��XeTh-#?�ʣxd.E���$VF'��Z�F���qY)�c�5�+dF�wH˘�D�^mѺ7�^]���r���8�sjr���6���6"�d c׏����˺��y�DԹh;���I%�ݬ)��C�(CP��M�3��pتe�O�R�Y3��I����3TǍ�LSݱ��(FY�ڮ��`̝��~aE���u�2� =��U�?�ek���r��2>����H���A4�Z5`�n�8������Q�E��<(��>q*�{�b������ �bBY�(�B?�(#^i���	�?0T��U⭊�/��;FB���ac~�!<ԎKt��RI������`���b��1�0UYCstsL��8:�$
��
e_c%�GB�3KM��:$����� ��Xn7�Um�o_��x2�[i,�t�O���GC�ښ$�+�d��}w}r���"�8�vк�?�P*�+fZ#�2p(���2�K�%��ڐ��b+�}x�������c x��W�`�66O7L��x���x���0�2�p������="l�7A�w�ǻ��}z��|D�Q9G�6�xm�
�o�%ŵ�V���P0���A�Z��`,���<`�0f�I�b�=�J��}�|y��L����-b�`;�*o��ͽ�<�w �{z=Mw���b���|spv��r�8u���p����7.>�����>�-�=�� ��wQ��ԇ�-Ȇ"0`mڷ˫���4�F'&����b�vƑu~�QF�S�1͟�܇����n�F �u�rzOR����k�y�D��;����w����8Ov,+3�;�3�Q�TB�;^�~^E�d7S��ĕtt7j�$��_`�R��6���>������ F�3����ݢR�$����4�*KH-���}!���j�MF;�;D�#rHz�Ծ��lr��T�����Nإ��"�V�>6��1�}׭)�O��/���N0D+"��N�������zz������o(��anΰعc��] 3ZI�<�+W;,�Y��zm�WSuݲ�mu΃z�KbM��?B�f���Tl�ET�V�~���+y�os2��{�*g�M�%!T�t�����围�qW�_Y�GT�|E�#�\��+ˣ""k?QvZ"�s�H7&��&qD�����:�U��&����k���e��4��FQ�7�io(�T�l��K����Rof�, :3&�r�{���kpT���ٞ�ƫ*�����[�kr�f��Bi�փ�z�����N��8���W`4��D*-Y�
,�0i�s�4����4�9Ύ��ka��w���~��I�]�E$_ss�h,ħS�d��鼠���I"��P�$"67����(���Zt�ڵ�:�ي� ]a�i��R������>�61RB�W�N�*3ײ�6�ʥ�@=!7Y�~�[���g��ĵ�Ra�3�7����o�A;�����䖍 'r� ����O�Ŭ�
4X���"���{� ��_�G��Qa�"�
�w�-P3RX�c�K�R�Cz��iѱo�ߕ��v3݊1���"xNr{��m-�����/n���[P����]��� NkE4f27L2m�sx`h��;����+�+�?t����~uf���h�Ւܭ���r�+�L�� o�[΃����}`���C%�D��P�� �Uʹ�8�ݮ�>��RQ���P���k�Wts^��/�[q�ĽF�ܨ��ET-oǇ�R.^�s3P <��;�4�㥅�a+Ȋ�����)z��M�we�����OU�������a�ˁ�����/4-�����q	�u�ĞN礳f�:,���G쐳�ɬ��ebe���8�8]��UPGA>��ѽ��#hl��S��\�n���Y \�]��m�Rb��i�C�30�� �1�P8z�8v�&��:����^�:p��o��6`�O���(�u���;��#g��A���$_ڶ|�=�c��ו����9��NM:�/s[��:���#-��~P�p�������z���$rŎ��{�G��䕧�Y$�$8���ɤ��@3������hG��ͣ�º&~1p��0yA�<�W˔���Zd� ���
�P���,���ͬ��/�����p�-���J���%oj&��'~xW��^U�f�Hj��u���+ɊY"�!��ST�PT@���|�%�-�ng���4��Q�8�G�Y��e��qR!�N't�)W�O$f�&b�c���@}\-�+FK�����n�xn�f����%�Qpلv'm�ޑL�d1�t�~�_��"	%�	n򝮑p�Y4x��}D��1�`v�y�%P�y�N�Ύ2���^��ԣ=�e���fq*��8;��sJ-k�J�ݵO�(�#	a���fZ����y��|6�s���C��l��*�j1f�ӟ��L8�,Z���	�X�ߎa�G֐lY��~�Yu��C���ȵD��54	� B�[�U4�����M�,^�!��l��bR�P)
����|V�af�Yam�0*�ٞ0���Ғ�!25����Ayb0��٩��#8�+��<?Y�o�-<�۰A�ݬ���)��\__�}<�`Ħ@��JR/v���c|�g
�?Ɨ���;������_U_�S[*-�B�����	�������,m���R�9k9Y�!d,����)��b~0�0�(%��,B�o�\�n7���U���;P��,�$x:}%U�Aal U����� 	������o�Jg��_y�t����g�K��:���帏�;T2I������{t�O�_��9L�g�	�w館�khF��� ��}9]�R����'f��8�B�2Z��;=Xp���%4JL�d��/1k�Cf���Ȣ�?�Ox�l�N�hS��N���G@�?v;���1b���Y���7r��wc<h�i!�GdF�$��K���p��z ����9멬z�D�щF`��jea���h$��E�t,�J:%�0o��>M�Y�����eܱd�P�5c�V��l�z0BbjrIk���
H�����J��;�O
[�^kT<gn��F)�s���2K�r�����AO57ɒz�EiԚaa;��8�ᘐ�;@��;�V�zr/z"�I���n���hi�ξ~���'���.5Fk��Jq6Lܚ ��9J��-�J����� ಾY���8��r#WxV�?���@�7Ε�C�����1�Z(٢�҂(���.*��:Rʑ�A�.2?�ٻ�u���3�q�@�� &�s�{�9CQ��/��K��()�ou�8<
҃[/���hq��15�D+�T2 
��˂��^�u�Gk[����U�u�3��e��ǜ���*�w���-0_7�F�t� ~�q����Ӽ�\+?�N/Q�?��	�ʂEcg��&�.���5�v�[
C�_���2/��� >�s��Fb��!t�%� (��ٱ�(�>��<��"�!vE�1΢���=���>OP�Y}b�D�S��!gE7¸�9�t�zUh��@��IXѦэ���-cH]I�9�/��1�!�K�3J�����懎	�Ù������^-�f�q���M{�j!@��)I�p��Q���7����<_�Cs(���%[���z+ �hY��+��5��ѯJ��~lPD+�6�<p��,�/'9��ח�->"�	���W���Q"!*�Ui�l{��b�|��Ml�.�)�|}���N����X��fbz��k�\>U�g=���8��6�O�GH���L��/ؠ���94��lI�J��0���}�_���� ���@:��?���K&��p$��잓6�2RD?��P�@�U��hk�i5=�uy��w,5�.���+����6%��|��NxK�ౡ&/4�,��D����h��:J�C�i�R"((��E�'������Ә��ʹh��,_����H�B������Q���h�����^(���O@�x�Q? �N��\K�ě��;�W.��?���6W��F�
fB� 5��#6|[��7�3КЅ�#��5��.���Wͮ�U�Ȟ�NCȳ�F���ifd�������X_%ϓ����)uEǨ�/]��slhs)m���
�$�d*�� � HK�������DhXp�������8j�����G���r���ۃ��e���0:�������WY��D�F!�FJ��������L@>��<��vqe9���L�/n[�8�i5ϖ�?�n�{��;wXZ�j$$��TJqn�z
�����/$���ɫ�����1��[�sb�t����*d{t_�	�?�`$2oj�_�����,(���j��)W�v���-��KeǤ�F!H�i����;x��X�es<�N��p���F7����{���hRJ�K�f��9sq��S�{��@r�n]�6���6��u̕	�A�|��F[S��@�Ż��^k�?*���'�E��D)�y���o�o��ST��U+�E��u��M,�'$sO0���%W�|s�(���^�����o��1��36o
��MW���#�����D��@wwv�Ȣ͜s_;��X�d�\��ܮh��5�У�Էo��}M���O�&�k���f�A��X�$&�U�Ym�:��rd/�O�~i9X���6�WI$�Ӛ�P�j"|�2]�V5�k�촚����꡷6lP����LS �H ��?��l��(�"�-��_�' wM��ДA�I��i�&�j��0�3#��14�	�8�n��v�i�0!�a���}�ɈsL֒�OW�:��<%Ix}f�[���h�`����Ḭ̆�����<Qy�tw�Y5������pQ�q��+�/�g��L�w�<N�BӪ�W[�:o���럴_7>�[T>@�H���y@�wN���^H���p���Y��\�]�����/���6%�>(^��S�L�g��'��K������&�H��tٜϓ�j?dUh�H3/#$b�J��iv!��;S5���=.=��n��*��f� 2�E$�ps&�k�-`7����,��,��*mc�	��æ�
	����!Q�ߌ�3Ik���Y��u���<G9A���閈�U��	3�lP�:l����Y��`3�
�qj�b��N��'y�G=��UA�d=6j5��V7�}hj����u���P��XCw�?\�J�E������8z����I�Ӎy��t��ߎrT�Gc�� ��J2uxr�(�^^�����q��|z��e�$�i��U{��z��X}���7V��u�5�n4�H����9��@v�D���jz�	
�|cc&n4,pe|aD��/p�CPl�Z�s����8��A�qz׏���E���~1��2�d�!~��{��sk#�|#�pZz�vs���BQ���UnR�v�Y�����������\��x?�Ϙ�ZY� 9�!�e2S��n]Qx�ݜ3��I5C��!���}V�g�#9ґC3M���1�}��D�.e��Ɩ����ub�}����l1p�"���ug�T��}�����v1�8QpX��BQZ�ڦ����t�����*q�t�������n |{gņ�4YG �YH�ӈ���� ���v@09���s}i��Ў���ᱩj�ð�K���.KB����sx�G��=1�4=��!Ⱦ�+�t����W	�b��$� zN��߇�G�լy�?�#��v�:��"���A��j�����4�a�v��
���l�A��%Ӓ�M]��=|�d4��������"�v��QgMĿ��/&���[�&6��i�hH���;�t	Ja�v����B�M�N״r0Zlu�!%9�:a>�$;�ټ}1��{	25��Ldڈek��'���_"�?��U�E�I��[����@
��<�%���KU���@w@���E�aQ���3vT��[��9��<(�U���婢���:&FǂY!�c�~����8��7��2���j�	��\��#�r��>^�����$t`F|~ ��7��=�1�E�L�%"�����g�ɠC�["�U/?�2օ�$�ڦZ$VD�:��[׸��pv0�$V���}9�{��hV��DWK�{v!Z*��D�������^���
����
��g<��y�8���r!8 �J'��"e�Jb�!��-�0����n��ph��?��z�C��a��~�ou��]�Q/���Nit�F����ָ�w�l]����mƅ곕*��!����{���;^���Q�!"�2�}�x�p��]��dt���M�]"@W�>=��W�k�D����:��KzC��[�ǹ��P����U��H�zWu[7��s��V����bQFb�}�;�-X��e���:����]Tq��q��Ƥ|�f�՛Ȕ<aU�/��p����t; �e�D��=�h��O�Ã�Y�U촤E�>�Kk>(s0�6��h�!S�"*�"����#?��5��"�?�xg����ث�!�U�"��]q?{��Gi8a1@�c� T|ne�SOZ�3�b�w[�<	�%��՞��A�V�R��:5����ۻz�&���<��}9p��	o��7CO~P�p�K����m���a?�?��e�1�=��=�S��ya��g�c��N)�B�=�|kX�K����Ō����b8�{�:J z����ư�3�rx��`o��������<�2�����Kzuq�UЍ�)4�Xt�u�����ו�Z�8S�Y\7UHP,Y-,z"�ZҘ�+L9{�_x�3"������"���|���q�&}��s�����9U3cѾ�3�m$l1��	ސ��F�m���,j��������Z8��Z�9�l�~�H:��ڒ����/���=�RN3zs�\��@r����QQ_�<Q�
EU�����x���p�=	&��7r'��;�RM�!�)�1BZ��W����"�.��#ű��༿!|,^�� c_�����9܋RȨ3!�4�\��i NI�b�L�y�"�r�z�����" /�Q�ެ);E�|I��YC!>��n_@�z8���?����΋ˠ���q>�z>H���&�E���	U��/�dpoe���)��O~ v�H���6-.�̮�5�E��L6&��f{��"D��%���-�s�;��0��Tk�ԡ���{�V�����z��O9"Ơ�w#�P��N�LZ k��ul������� %� D���q*��`k�W�̓�-�TqvL���s1��z���2���������jI���۾v��<^�P��Ȼ��M�.�V]���ɬ2�_�WD}���o�,��^�+-�����]���ZԺc�k)��5�� �y8fqËd�}�hzb�ݗ�Df���S�Q�"�����)lv�t#����3(��y�D�	��Y�'�i#$������.۲b�����&T�)<��J�0�q�U��>��p������lǻ�������Y����j6z�h����N�{����"�Z\�#�7�4��40(.˕g�{d�b��H�DB�sm8R���0wg���>��i|1YD)��Ӥ�"����<���װ�r�}-��M��nY*�J�s�_�u�NU5o���x�������N�kq��*R���S��9C2P�����eQ��;ͧ)��l�1=�� K��'Q[{�t��3�=Jў���������"-��*�*s�B6gR؆�`�~�����|w(�\��n�?T})"���e��ǽ0(m�p,���o�(V�|�1�/ׯ�ڌ�ŠTw\��q�^:�i 7�dcEhזe���يc�!���4t�����k��o�^��u!OA�v ��ϵg?j/8��	�<5��`��z���f~}��v��KJн���v9u�w�H���r=�^=}��h�f�ga�?�k���o�"��<E�-�Ґo�+�s�?�ae.͢>�|.>c��>y�'� k㡛,��I��-�yP󤙾��ː����f��Y�i��E��<��}�V*�1,������5N.LT��FU�-��N�/G��c��	3��CF׽�.sڸ-��}��)OsD����>�RѸx:�����f�v���f�H���nR����v��Zd�b�Ɂ��))L�d.s���uDu#��ƽ�\̵ ����iF1Ù�}pr~�A��^��S�w[{F'-t�b	4�f8� ���K�헡�|9�v�TOJDE��}��&����f"��\\�\�gY�fQ�@�wk��{#@��,;�Y�?�����k']Q'EM�sX(�r�Sg~��v\!w���{v �w2�{*�)ݒm[J9�YK!=0�\U���s��ܪv��ݏ&���?)驻>�����#a�S�G2py���6-��z;T9^͏�
(�j����Mxģݤ	y��������*���s����+rJy"�C��A�ݦM`��#νӐ7UFG��[�|��V��)��/�{��qD��4�[�8��9*u�P<��������72�o����;vu�ōG�c��'(���pK�W��asX�T{0/��w�m4I�����^9!��O��xw(4�~j��[�H��t
pQW!��39��Ԟ!�ar�}�y���>�ш[G�K_́h��c����X�B�l�_�!;�-�A�g=��<�;wx�x��;����P� �wa(tѳ(���i%r������ʻ �:���[E��J;͓q}0��_h�jמ�g���S9���}kN���rf�7H���N�(�X�'M��M�zL�Վ��+qE����j~a�h�UŦ~)����j���n�k�@�RQm�`�BZ�y�=hS�G �$i$�1sl�/ a.^!{�5��U"shD�	�2SpQ���umB
I���}��UK��T^#pv<���I���<G,���1I$� HL�����������<M�Q
̆��H!�0� j:�B��j�G5=���va��@VX���H#�+�gW^��&p�	���s3XŌ4Ns�[t��*'Gʺ��_Ί�qXQ���X fu����R�V���� +�hR3b�*�1^��@�p��N4��1�P�4CE���ӷz7Vp.���/-�m��Ҩމ�����g��	RP���[���{�gʸo�D�{�6{h����c<y��hz#{ ���	7dDY��ۖ�N��!/f��a�el
 3�=�ڎ��G]X��VkL��4!�"��ۅJ"�-�^d��;?��QPy7�������.*�d�������q~9+�6�-�y'�0c�?�EK��ms�2Uaud�}&]Lz��*gCV9���|z���ݤ�l�y�7`�_�L����]���4�(bm��%R�]��j`,��=��'r�0��Y��+��q����`�n�q�w!�H��y�d���c�\����U4���j?��S�#��)���#Sn�j[�k�q�s��]�BY��'��ްJ����4Đ���o@� �U�ͦ�r�!�ա�ٷ���󾅋����7����
�o	~�X:�i�¥�ܞ1�* ~�֊@H\Pt����Y c���E���2���s�������jh������So�!�~^&{^/s���Qݔ�"����0�ۯi�ɉ�#gr ���m5�Q����O
v�(%���XbwFlq�UX�������lɺ�i�Z��~�fڀK��Z��ݖ?��'��p2�m���R�l��G���W.סT��T��B��,��F��cDc���G������Τ��W��:7N�����s�����k���RnA-��1:�	�_�z}���QFzNa�@�2W�:H�	_JΦ�ز�ESù��:������w,�A3qf�r(@��nLг��4G�Xh�3��>����B� |ټȳ3�'�*n�������u��J�!=���-��=��:!4I����4Yu��ho�tse_`b��Q��>���ټU�s�����φ�M�L�WH7��"2f��O�����?��� ��r9�W�����P%���Dc���p�#��r�5�9#N2��=ٻ��D/}�KP�4肯�nL(S��W�� /�v��g"NL�J
����|���;�,*=.a!�������TN����~4+�~���թ�=�E��7���ͯ��,�X>˄�N�v�Ý�=��N�^��?ı��K��z��l�L�5�E�;���/1)_�V`y�>�s(A�[>�Y���cأ��Ƅ*O�Sm�&�e�N����mxo�Zgll�q⧵L���u�-y::�?w@<��������/�M��'�ٌ�&
�ԫh��BWƝ-��K�8��BCF��uּ�����3�h�+v��~�"T��ұ�>ߙҬ�H�v����g�<@*lo����	L�x�]j�*�V��1	n�pb�0�v��~`�� �.��}�5?8���I�Y�	��KS⟊���v�~���=GmN�D�'����z�ڙ��`t�t�F�;(ۍ���*6l�g��)E�B��{;6/�'!�Ak���l�a _��D�`7S�u��\�UwR�O����S�����W_r��OH���aN�jl�:?��=9�vC��41�z�ޮ�r��������+����j��S`u��Q�DD�G�~�X� ��0�(����������Ԩ�3�`H�H��ݔ���"��q���4h��Fu@Zշ�P3Khb����.���$� �\�i0P�R7ַ��t�O�G��f�uB l/���6���b>)�]7�3�*��VD�d�Ћ���s���-J�v�����w�����{f�WǠ����
9u���
��pU�t����,l��ߗV�V�9�T%����t�}�j��ϗrj��]]?9�Q���u�N'��^H�{����X4�n��fs�O��65��X|�f�,�Gb�a:�K%��>�7��!��� ��J�d�4`�ۧ�}wT?��s��u]��,v<$�pd=m?c���l`��q;������d�s�H��07^mr<E���4��m��_N�S�!(@2MA�S���:c*0lr�������U+![��
}_k-��5��I��8ށ$��<\\p?\�S��x�M��OˮKJI9�6_@�Pk��<��eRekK0�':T��[��v��7��N���hQ��̿S���')������U�<_������XS��C�3�ڏ)�1����e�+t�)MM/��֪;ǾOfq��a�Ы�ACIy@�'U(����˹�JNak|~G��tj�̊\��.嘔([�z��贄���9"��_!7��1o�\K��%;��m��eyKd��?3�qI�9��Az�ܽgD"V�����;��G�7��N8��`�������mC��ى���D�3,��=�nc��ؚ��3��m:��o���ư��QB<}1ܗ��/.��o �܉P�8��-�Q��9��Zy[SrC�1�:\hq끫Һ��; �""o����s���kz�~�M`Zē���z�0z�H�5G�I�̚9}��W-O]J�(ڔ�K��%u?�hc�j��Z���W�{^\z�v��<�$�!C-�D>���T\�,�z�z[ߛش2�#./���!���L���oXN���/0-�����h%��<�ƕ���R@r�U��1���D�{���c71�dwWE�`Z�3^�<	����Г�8��6� �7FБ�h��p�5 ����y��a�G�$��h����W��߰�K��oBaS�In��1�E��1^��� ��6i�޲�G��"g��g�N�Lx�Ϝ|�]��S�
����dT��f|%���J��s-;�	����7�S�EO��-�.��i�@���a��r"�X�<���
<)���;Ok&uCpQ�|ӯ��:Q��c���~c�к��3$8���g�4] ��� ����M!@+��ng���˩B��5T��$�4��YN��Y�8hq��t;؞0��'��x�$�le�K
c��=ɺ$ը��H��G��C2(��C�@��v~c�Ĭ�;�]p�Z� :�5r�@��sl�p�ALL�����f�i睻7�7�����+d��z�-`��hJW4Ke�Ϳ6��>��n���cz���l��MKI�7��@��w��ϮL�(����t�*8��43�жwvxw��+�!��M�{5��B {H�>ů���?k�T~Pǩv!�R#�-��KUu�t��K�)̠��7Bfd)�|��E�_Xˉ;8|��{a�������W^Z%:w�|�O�yq7�*�yCs�X����h(��:�c����V�7�M|m��;(w^؀I���	�ׁN�5��^��DflS@U0��b��}p����1N���{�k���������%pBsďr�b�{�w�N�L�i�z�c����h|���G=�e�P�xĎٌrz΍a�����`�"9ۈ���xG�/�� �L�n�I��nL2������E�u�v��z	He�ʏ�˭N�Q�uJ�=������_�tI&��ح{���rHf�E�-����~V����|J����	��|rԩ]3�E��RЈWo����S1�����K��H����~�aG�c�� .�:���”��'˰zF �+H8��p/ �I���f��>Sg ͮ����!NZ�f�
�DJ���+��z���4�q�܉�@VI�#��uհ���fb��G*F/�?�)	iV����6�C�<'�/ n�I<W��k���P�C`�L�!�����>D���4DZV!��.
/���c�u�qn�e���u��;��`��?�^�C�Uk6�G7��\���e�9l�� �C�BL�#����ˮ�-=6��	������w5�ٟ�,�v���W�9�g��[6T־�
�<�ܥ�~'ʄB�0N�!T ���5��\!/�ˏJ�s��^kE��;�E��Vo}8,��#΃)���p4n�P�뤺�:�!ڬ������6��ўP�i�u�+Ý})��i ��®��G&`�����TL�^RwA�ce���$7r�A �+���z+m�C�>v���Y���D�k�	��NӋi�jW��Q���e���<�W���{��(1�/�6	q��Ț�v9-R�� �°�$��G=���ȴkS(%��d���i�R�A��2O�
h��_�([��Mb0ҝ�?|{�ٵO�h��C�iտ��10��GW�̨�và��VoZ�菪���5)������'K�+ʊ�@���!x�����SZ+�'���+W�Xv�M%�Nɇ���:l�
&V�(����=m�xˆ���T����\���@�?"4s�f�[��C-��2Z<ߟa8�����B���ܛgC[��|���um �z����-��.s�������U��$�!���-�X,�p�= �{�HH�t<4u��ě���̇��d���oM��e�D���Ҝ�'T�ֱـ�zX�`2�Y�_vb�)/�g�FpxrH<�[����ZUzewV^o�r"�5r�j�t0w�Q�h~��w�� tqSW�v+�-�^L����6�� �_�����
.�E�YY��?P����r ��c����+��]c���m��l��|o��;8�'��,���n)$k3�s��9	n��]A�a���
-E���&�(I1�>N6õ5)izO���7�EH�RXX�z��F�K�ze��3 >f�:g��	���&�'B���Hu�s�Ɵ�P�Z̄��*�{f�=����YTO���"v�_���5���8��0p�\Z�[Eו��u�[J��{R��qa4��xGe#g��V	R�C�3�f�/:@����x�v�J�A�A�Ǌ,�u��8�r��wQ���c�Z8�X��p׷�<������$y��K�'�-��,����\TT�\��J�[����hC˵��V�,���)֢�
�`��BD��J�|�p��6�����sk�x�ql�V^q'RHx�&��>��]�P��/.�Kb��19_�����+����k"SmN{Z�:si����Ma��ya�I��c,�I�}������B��#U-_�`�&AI�$�n�1���<����}�Fz����m6'����gB��'���.�W��U�Ky����>Gӄ|��A1ǅ�-�GB��>{����D����@��z�rH-M$��١���·Bʸ|ɩ�7i�����]����d�A�`UC�p���f-B��ٕlﾷ����2Zk�u�/�Iϴ�nkR�����L"�����9�Y0�Jg@�"NS�O?��+�@B	q��p���7�����Q�)L��?��Vq�4�>Ppp�0\�7e��h�2�.�����i�7#q�i���S�7~pCѢV�8���^��^�,x��� !�Y�N¾ǎ�gU9*��(�T�R�����y�7�<Ao���]��5�Y��iv��s��c�ͨ�*��d�Gy��Ⱦ�^o�<�}�o7�<�-I���U�1Oj����x)	��1��H��J+=�/���}�"�����ma�-�����/3ۛ�٭��^�gG�j���s���'�7��
s�JU|�8��"x��;�bi�.��T"�u\ ,�f1����9g���ED7a����Q�#}B���q�V�)��fj!+hK2�U��nh�-E����� �x��w�	y��(*[��;my�%�����JI;�贪e�c��\�F���!q�������g|$H�Цa�K����Y�%	XW� ��I��bE�2,B+J��u{c*MvAM�IJAj�Vl�>c����(x@�ak/��nJ�g�8`G���vF��"*���.'�`B��+#��_)k x~y�������y�`\
���se������V�F�q ��Q�Iy��G���Ұ7;�D��b�Y_�I8�@�V�2Pט�g���_|ک�(����5;��p��d�S��t������ �K�U�@�a	�N���fj@drL�G �������p��$���[�=�!r ��]��� >�_ѹ�}�X��pwtM�*���q����2!L�&&��w�����}��od 7�k��1T#c֨o{��n���	����ثƀ�^�ɍ�{�r�{�Y,A�����z�R؜d������ʪ���&*2��yRɇ�h�D6yi�t6oھ��g�N�%�5�yvc�j/�j��]�'xyH45�G�6l�����en� �;5�zk���\�E0�� ��L����$���D呓+�%[�~��EcQЅ�'ҳ:��c�A�382B�0n����l;�W��L�
���
Ct�v%�2�?iREp�r�z'���Y��o� B��й1%�D:�F���b�"����6�.+ݙDy'���[M��Y[J
} "!�(+E$�S�œ������2Xf�N���`���*w�A�-K��ORk�\-m�eL$_���$�t���6���s4k�� 'e�4w��%�Fg]<���"��mu��	�0m}#��j[�C�����k�Hy� '�LӖ�<�,GԒ[��3����:��6�Uu�BӺ�L�n�8��e�n��n�<���qI5�אq���Z_��@�M^y+�S�
��8�(7��- �ak�f��LϬ�8>}�X��#�5��I�4)=��#�32s����+�~>�6#�s���eē�i����+�ao*]�����G1<��	�#���m@��\�@��u0��p���p^}�i���o��aA@��:�p�0�'i�j�p�Ѷs��5��@X�=^�p�Y�3�H�#�r��*+�*zf����SC���Cw�6P����H�t��F+v?�`� [9N����! ��P�t�'eO+��ȉ�2�3��v�'43n:����%ΟnE�R	���h�^^|]f9��S��e���d�J�(2�Z�D�J5D� �y���E+�#7���p�+�c�;H!9����#�c�A
�g�x�̷!\�ǽG�rx
CƝ+Z5��AD���e5(ƝA:�'���z'���e7��xQ7�5)}S��d:a�Ϳ~&�����0l@�D"�;FޝF���\?i!�"�D��d2F�y�%y�Hѩo4��0�=t̩�P��X�bw�խ�_SW6K���SN�aIu�;V`K,.�C	�����9�`[��3�訠I;��^�u8�q��ޚ�x����F�І�)�q�d ����Ws����N㲈V��M�7��ox(�~G�AO���?ST��$ϰHx3g������"[���\�PF"|v����D)�i�Y~"��
��D�51�v��q�s�b�a5Ѷ�|��I�)?�M�诮��iAbْ���kL��r4�0\F�������y�V�V��X�A*rP�bY��T%eʰL�sؠ$'{6��L;���?-ma�����W�*޾�n����hi�ҽ�
�#G�HBtd
�v�-mz��*�'�|u<�G{.��#.E����`�->z+�*`i�P� 7�[0s�:�t�]����#.(�}��<� {Y&a��^��1ԝ��0M�^b"�8�1N×C��Y��M�����.S��]��n�7��^v��k�Kɳi�f?D>��Z�? S��Co�u�Y��<5��U�+`s�#�
��RQԛ98[��%`�ϯ*��y̖�����\�*���49��D�|���K�z�^8<Q��F�(j]�cf������>��S�'%�\&�T�I���.42�3�z��x��`���
F����p[��	��� ´��-o'�
B�K�����eZ�V
Y?~�b���$�Y���J7��"�ai%����gU�<"���E��Λ�:�fɦp�='�^\Ӱ�;$�-��/6��ht����B�Ta5(���A޽�\����nn�G���9|cKi�AM~<)�[��'ȃ�՜�l��]z�+��v>t�r%
jC��[�j�%��:����3��(^S�� �]H�;`��*7���"��6�t�ϓ�EI�4;�p�P ��_V��g���g�"��mӔS�\�	ii�f�2������+`R����,(_6����׳�ͥBr8�d`lEu��C+}Í�C�xf���3���UA������ܢ���"��DY4�K��S�X	,�2h9���LD��`���r�r*ȏ|F���|����7D�~��l�������|H��h��,n���/�^=��Ei��I�l�w!�Vl��ak��g;��	S(r(�&y�[�a��/n'��U�/h?Q��;N�C�G�y�U5������ۑ2�@�[����I���۲O�۩������Cܾ'�
�f����ipY�U�Q��2h4�DxLÁ%`�r�-kF�=��� ~��d��r����̲c!DC7�Sa�J?�\�E�(�]�k�o$������k�/��=��*�C�I��S�{�d㍖*Cd��{ӟ6� �i �!�C�����k��&�}���Gan������ jY�z������i�\�d��Y~q7
��n�m��l�")s�!.5S�n�i��L�[�&EE3B��xE�*x���`RYD�� T/��Pt$��uWhU{yrҁ���=z<�N���9�(�G4o�/�A/�1@Ze����U�Cֈ�|`0Φ��
 /[C��So�"s�u!�Ms@5R66  ~��[�1�-�0uM��[�K�6)W�_*0�0����Dn/�
[g��GF�qUa-�	�΍��j�A�n3lm�ʥ;x.�H��g�/����_~�sqq���	�?��뫐�kq�=O�@�BC�D���%b��̜����V����t.n��q��N�}�wP��G#RC@�X�=���ȟ�4`g�6���&Q`Ow91Pi�Nu�WE�*���`�b�M�0Z�n^�m�÷k>�R�{�n�$s?��K�,]!ˡ.�"����r���J��^@[��J��������g��d���j�l.7#�0?mޒ�rڷ��P1���S�G���
tL��)���1�7��>�����8x�X�0bXߙ�R�2̨ت_k�r#��ޯ w�<�P�`<,��`��B0
�JR9��חt"����;�����x�b��]�*��,�?�d��ա�gߔ�#0�u:Gx`�XY�=���e ZS�+c�ŋ�]�S��:�� ZS�����l�X�^���������*�O�����ҹ(�k��aa�����b�$��Yw�<v�%�֡o��-4M�K�f�5C�A�-��t�Eo�W3l��|O�]lW�l����_��Ȧ��j)XU)w�E8���e^,� �<�k�J�z ٖ �>�WIM��+r��>>��p��Z�.�g�`�s�ié�ͭ@p�k��>�/���xB%cnX���
]D�yo��3H���V J��D����.o[Fh-FNb�E�IkS�?��7���ݭ��MM!���;$|z�BI?��Nh��Տ�y�OT�!�Ǘ��'С;ZQAWuת��.4�`"^�]{�u�mݟ��
K:#��<� �U�7yb�F��)�~ړ�Q��5Y��+���'���_E����f�kq�ٳ:r�/d��"j2��&��(�v�ƆOC/�Slr� ��ܢ�҄Y9uą�F'd^�f�6v�D�+{:��L�\��s�?:h2�����u�p�����2�lMi��A{�v0&����P���N���L
q2C5�O=��ђ6�x����v"�׌���U2��1�_7�W
��k�(�s72�	5�?�����X�Rq���;�5�9���[K���+����ÂƩE:���۽�oF���Xp@�p�j<�4в	+E��L�y~4ڐ�{�C.]c��Bso����Ӡ�9n�����L�S��V|Hz9���Z�1���{�F�-	q��E�7�5Y!�0������R�)���uʲjU�*��j����h��R��ɮ��n~���kJ���JΕ<bq�l/�5p�V�T�h�c ֮}
T0�j��~F�#�F�f,:.s��U����J����&հT`��d�#���Z_�����&fp W��V.w�6���"�s��%Xk�չ��3!�=O�Hc��!(p��,�>���t3������7e���&���c��V`U�X�4H P�$b��o����[O"P a*8�3�� �uJ�?�r4��Z���2��KD9�/�-M[l ��9�t�@�~�Tm*�bHjVK��ΧA񂍽�j!��ɀ�v�&]�^�s7ZI�14����r��k*_>?4-e���ө�Nf�[$/�{�XK�ιu�k�C�(g,�7�͋�GI�eLt��*K��?�_n*ۈ��f1hф=��"��r�C������pЉ�u\�V�ӽ�;*��>���F�]���s������8��.-����A�j �{6y'o�x�:�(���j���%t��L�a�R�P?�lߢ�zF���Pޜ��ΰ
��d���fv��f�
.��˂�eM-%a�M�����.|L��-�\ d�}�1ϓ���#�ڱ�J`�i�)�<A�^v��T-[�B[޷V
��*�R�T���`�ߏ���������/�����b�x�(e 
)�ƌIZ��5g��1���q�Fɿ�N���P�W
T�`/�.k�{\N��s�{�q�$x�OI�c�mq�S��TJi�����������!�*Q� ��'��1�zp"�	D�~�Z/�FY[6 E� ^J����6�p�~P��z:��U �҆�M �n�?������f�,���f�J/�"��0:|�O�:�H>qʦM	��Tw<�j=�tI2���Ԛ�{�U<[d`g�����[��W��&ٛL��i�ƶ��w-�P����G+=)$H0��R5:���u��l�߁+�Ei�d�ۛ�kWc�X�M��	����)J*6���y͆"�l�&+�h_���e5(��r�}�R�jij�������)��Uh���)#����T_z�8e��3�S%�_���V9��nV�-.Z�����r=
���Lt�vKM ���s�g���6��.g[�z
�tڗ|��sM�y�N��!5��mRm��J��.�0�]2d��Cp\(ʹ���!��m;�+�Y�T
U�6D��M�ד���z�d��[�^�G.�� ���in��d����:譈8��'P����>L_᢬��U�f?ꤪ���I��<[��aO�!4��. �9L���S�B7�FD�վ��B�B�R����P�����]��G�]n��'���Z���v�/��X�MQm�U�Ηˎ9/�H����u��la�/�{�L����Eh+N� �/5�B
���|'Zq���B9�`�f��7�|�{�C�e�`�R�
�5�H�~��a���	v�b4���*j^��[��KU7��hE��~@�e�^��-Oނ8	��$gI*+��j�_�@����@���C'p����d6T�w�5
�̲J�7����Q �]�>z�Ie��n�+g��S>Dz����z����r)ߴLI�O(���� ��C$đ-j�2���[d��z�V�da��\��v;)�#I��s���'�k�]����˥��$��#���+PB8����8�S~&9C�,�Z-݂Qd�G���Q�j*�� *OX�D���S�(XIb7�#�㕘Z ��_��D$j&N�y"�N�X���#�L��I0d���~F4)��t	~��U���KKi��7�Jx���\��jq������5�����^��j����Ȣ/#4�Y��'1�l�I+�J��&�BRD /s\�u6�bIQ��2�v٧u��u���ÕNH���-�x�����S��A>�B�!N��h�i�\cnI�����M�׊�h����L��'u>!�F�u8�0wu}���L'w��)��f��VW�@S�uK!�R��S��"Ν��K;˅w�=ȷ�c�|+v$T�cݺ�p�luq�E�e&g��Ç�0��=�N���zdHLM�G�7���*h�^��!ѽY!�s��G:�VFij�u>+���X���_�"9��ɊE��y����p�5��0X���7l'�~�X�B����i;|̫lC�YiF�ZI�
v�޽� Џ�^�&��Zv�i^�(��y�uD��g��Ǉ���(3��[V�OwG�(�JM���3	Hp -V@A<�l�u�,u�+U�� ⮹JT���u��>�;e��Y&|f&]�"�c�3z�?����~lfnA�~��vm�9}�N���>�09�E�?��z��W���U0x��8D4	D:�g�7�����0�3��s\ƣ���:���\�2�2/�#8�Ɵ��P[���%9�U{��l%Й���lI�yC�h��j���'G�K�*I�:�8ZlB�:i_o�7�'M�l㜣��
�HA�����L�d�c��h�p�4Tȶx�����>�wӜ�*8�IY:�q�h傽<�:+�����d�Oh������_6b�H��놭Gj�|+1��}�LC�2����5U$��b�����6��X|�zX�
��t{P�;���~gL.�ڰ�'���|,5�-+4T�����[1�Ǣ�C|�8�Sq����ܐ�L���&G����'�� nu��w��&���Շ\jK�]o���������I���pt=�ʴ��NƷ��#h��fT�^��/6����o ���|%�\�<�'[���.3j#���P,�	u��;�asQ+w8����D���b��3=�XT�����Roeq������9���v�M�鄲���v�}��x3�(��3Su! �,UC�4�C��	ڨP�(]�Z3M����$+0��D�Y�D/�{1���݀R�s��BO�檝u ��=���f��{�WڠҔ�F[ܥl+@�I�Z^�7V0��d�@�x���wK�!�i}���Ǒ�1f��	!`7�ø4ȿ G�AdG�t��YO"L����T�8}<�b�Q	#�J�#���i�l ����M��dj��QD�\cc��zNׂ
D� n��/j���������p�C$�� ��8�X�4�� �.�ı
�ٮ�@�i�"���.�(u��3LA���2y_?Sp�3K��$�!X��d�kc��@'�=���^�1ё��z�a�~���%�Wǹ�\�q��=�e�}E�&��go�B���f
�s��n���~�+&R�x�]���V��jd����M]�Қ�  �x�k��[�Oۅ�O�QU\�&>q��pf�)�bP�fkΪ�0�$(W��X���H�����:\����kl�:o �W�L��c�d��J���V��:%3�R�����'Q2?K�@r���!I���k�b�1�M��A�'�2�c�Ǖ1����Kb��g��_ĵ�ҶpW<�1fR��=%tS�Wi(,�)�>)l�r�	�A���{8�l�Z������C����eki�
���&e�r�}�0T����X�+�-ݾ��t��Ț��F& m�QJ�MO*�3�&��
_�D�[k��Ee?S��1;�'�J�m�b8����xQ�� ��n�m��c����j�'�)��څ#��y�ٽ�dj�!�)0|�k��ֺE��k���{��v��(C�m#v60�t�yI�a|t���:S~%�����%��E����Μh��+�i���"�Ƞ>� �B��pՃ�~�ʨ��>0���Ϝ]A6ϛ�i�ٯ�v������^ϜMJK'@_'�w��)���J��R`�³�/Re�ު�q�OS�?S�&Y���ɄӒ܃�^Xi�B��`ٍ�Á��,(}/}>���W�~^���[k����Y�\y�|���-qQ�+v�'�$�/�|��fXB��xEqo������I�٥�,:yV�5�ZGG����K�8�N���tc��?a�Ʈ��in��9+:̙��'�fs�p��;*�CD,x�y�1<��f7<�!:�#�n�Y
�1^�8�i�~7��v&��ʧƷ?Z�`3��{B���TIe	9�点��\��u���̍��b��y�'C�?E���;�}�ǐm=�a
���9p��e%�aZ"�}���y�����p͉�m�ɇ����a�����X���-����«`�(��"�z~x[�z�ĕ8�1����+,d~mY��3���l�5=v{B�J�4�"l���l��<�{��@$��tp��ׁ7���A�~J@GZ}�@[�&�!x�g�Ϭ���&{��S�Q=��)�û:��lIǬ��qh0��1�(c�3�~�`+s��fxڒ�'5=+"R����Q��m]��LL��h�!��T�H��h\gEN��/cO	����g���:ᐺ:��Q4���Շ$ٳ�<���rm��/@�k@�Ѳxhp%7zR��x��ޓ_��/Hm;�hl�c��>���<{څ�f؜�tD�*�CU_��?����0�������ļ[f��v��	����$Q�֥�5��SL�(~?7��-,mej��ڊ5V��RRq��[�
���6B��L��B���_
�r�Du[��
�I�??րE��-��W:li�Wl�������,8�$Ae� �	\&��U���gh�U��ױ�܈P ��� =˳$����m���hHv�t.���M�3�.��äwK�(�w�T��h�C������[�NJS:$r�a�o���\n��m���o`��0ڋ葌��pC6���5���P�?��	(��������8a�% ��Jy�o���g&��͊�KzU��N�q4q��5�]	I�&$�!UטS�s0î���
�}7���f �,���ne?�4�>&���1���)�P~�h?f�ΰK�:)����`U,j&Z��(���g��0�0��L~n��ʨJkL6���i*���"����*I�f�m;�1��)Gڋ'�K�ឭ"��Fc����mk�MQ]��\k���g�FMNǧ��'�Ō�)�����J���K4��~~��8e��R�%�b���H�w!2�P �p�?�}�)[��q���S4i��}X;��/��b�a,XԴ��:	���`<�u �p��(I
#��tB}`?�B�@�.K6�y���WG/��Ĝc����� 0E�Y��Rx_�TW�����Q�O�m=%=����%�6$���S�k���A���zO��:_�E��%��L=�����ퟞ<D��uڸ)	E3F'N�v�ڒ��aɟ���&��J�!�B���μ 1��;K����R�d��Yc����A�w�5�d�����j����C(y�l��v)O27G�2�h1A���N������}��^I%�G�<Az�6�ͷ�W~š�Dfw�83�*��a\�~�;
NgҜN8Ջ]9m��L,���o`����F��4�vI�;�k��փֳ*��l/�,���c���5��z���.�i��S �Ŀ��B�ɴAv��z�E�y3��2�z�RvW$Ѩ�*�=�g�Tr��;[C'��0��*�K ��zV!'{x烎tCT�dU�X�(B�<)��.�Q�-���D��R�_��)���P,gk�o���F���?�ܝ;���3�Q�*;Q�ߑ���P�ExZH�?� n��HXt��#A;s����_�N�f	�3P �k-#��px���0;c̦�!�����G�Й����'6P�^˾�*��u��28"僥q�����[B�M-H�ۍ�3@b�"�|J~�Vl�SDL���\��bS_�vƲ�wOqэ��´LƘ�{�0/�s'P �/���b?f<t�x�tUZQA�Uieg:��>l[I"��؋{��x�	�d��8I����Ś>�ͩ*2Z�����r��`6�b��/vE��R$�߶n��x��d�����i��:���ȥ���`?fY�%oQ�M�$f�E@uQAO�m��k���5�`�	�il�$����rH��ht!�&�\�ȒՍ.b���{��WcW��o-�Ե������a�:�]�CX?����0�)p�<̎)֋��7���\0
j�@����W�eh�.>�*(|�A�	S-�I�u\��>7�/,)����޼j(� N��Tr��/�48�M�ʂ��Q����~b����9���}$��_U��<��Ȥ�� ����.z�K� F.�-��
�I���1���|W�x�(��ce��/�,���Խ�U~c ֜�C�Z}���[u�v{`!ڂ$�������#mA�j���z�?�rKH^��#G�N+�H=/�V�/��
���=ƽH�O���!�mr �[�l�s���'#җ��|I.�O������B��w���T0�v{��v`sV�dIC�� x�?����xk���Q�����af�fg���,1Q��C&�[���Z&u�+�G/J�G����<�ݺlк��~T-��;:֖�cP���Ň�Fp7���l��^`�_ b�T��<Wgd���U�㏫��	v3_ܔOS�t�c�v�uH�c�p�p
�U�m-l������OCj��f��������6�lr����6���Ӫ�t�hN���ne7�UK�Н��Pk�k�kK�欔��Ǿ�Z4x��!L�Լ��p_�E�����o�:�+zؿM|QPX���#�!R�g,����m@�0w����E6�kDUKL3��?}���m��۝.�ҫ�}��&�G�׮��jv#���@[�Sny���0`T�%1����qޥ�a@A����Ư.9�2\k�'�3x�2�����dr��G�.��*����A�e��$��0�Q����&��M�hgCV�h@d��7Y�>��`�����0���j��Xw�{�5t\bU"�>��fm�[���Q��|��(r�?B�U��"��ge �!��+O�?JW�Q�ZJ���q`Dê�uI,
�� ��j�?�;����l'3&o	�qQr��~i�.�����6��Tl~��� {�,���n�������)��k��Xs�e�.h��:!2�T%O���x���Z�B[�|~��9vi�MIs�؄�"��J���a�������wٔ�:��5z��z��n��	�\i"`�|�;�&)���᚛�s3|~�k.�l>)���١�~^Ԫ���+�?d�֎]��cU�w�贻��	�
x5JA���^>Ԁ����Sh�� Z�1��|E5��}�m��p��;��`d�l2;� C���M䱞M�j��n�k^M�w�;�2<�u��|�	x���
����<Qgj/)lu�j*��B�s�I�m�f��pI.��)��w�IW�c��v���2�-9�.7:���W�Z�F�?�����'y9�` Y���ၚ���Q�g�e�P휆�FJF-�v������'�>�lU�;Zp)�4�N"|��!�,IK��D5�;tE��W&u ��O��j�P,~%uC���Dk���I�f�yO����Q��7,�UyQi�܁��c3T_�q �U�f�n*!����BdY��[��7��bPҭ��l�\:����ķ�K�P�������	�=��~�2�'�6M#Q!����t8
��5���"��#8��	䉠cZ�Ex|L�s4M���й$���� d�Uu״$�1���͖�b�����%rΑ$9;^j W�WN��ܚ�Ft[���'�5�)F�1����ҟ�ˣ9'�b�A:��IwX��dxqǓ��3�2�t ���p�8]�X3�΂E�cSgg������9� Q-�������>��r�*-�OU�����hR�@��5?�}��_~?�]��}¿�ȳ�3�K�v�E�u�O׎Nt��n��ٌ0��姠�h$�<
�]�e�1P��q�����-~��+d�q57����8!�g3��/��]8�f9��� K��+�w���˚��/���	,���[�෶�N�0�0���W�xRf�/>;�n_
)bC��ע��%�Ҏ��1%tb��pXŤ��J���H�u>��(B�G>"9<�/��8�;e/��Q	�2 ~$"���rB���ѪA0����������e�{�bxQ�,�S/���|٤����"�T�M1D�.w�P�q>"S2��}eL�_��Tu-G�n��S��Ax=@e�(A~!w�k�IT8~oJ�i�	k ���"B;{��q�]-G>(L�v釜����ձ��[6�(*cF�b�<���)I��n����\�f=*��f�sG ��E����5Ǩ	0�Rϛ-�A�G5��?��	8	�ۃ��=�h��"��N�)߸{��r9�B�P{,���&r�(L5�[���G7 K�C�~�<7�b �N͕pv�r�y��Tq�yg���뜡¥P���k���������	��a��5 �{�%ᡜ�A���έoO��ɗ�ǰ�E�aJzC���)��د��o�%����ܞv]����5ɽ��{)���sS5��^փxk�� !�ɊQ����u������K|28�G.�6;_���4x��~']��l�*k�E� 
j�`"�a�<��������VFNډ5�`Ad�ة�K��N�0���b��������G�-�fp����;��c%&>��}!���_�f�cY�ʉ�1���������]G����	�q��O��i<��T ��6�֎����k��:�*�0!L��X�����ђ��`0r��L�I
�" ,'�'=�'3�����b�C��D-��`c8�='O�Pa���_q�m��U�E��䘩�Q�SN�#dj(3*���1+-<5�N�[G�Ǝ]'�P_��N�<V�~���%�9��O=ސ[�#��ց����0�\�ߗ1�	���9�[.��fC��W���8��@��K���L�a%��KT�i�����i�wƤu�Y-�|x%�#T�F�,-UQ���������i��D'ɥ����N��)Z1���i����JҲ_<�#eH<��;����v�1��y@E�?ߢ�3�X���!Yfx{
�
V�t���/An���X�QØ�h:��E�&��� ��k��Q�1����D��J�����~��B����Hr�s���@~n;W1JH]�[/O��MP,�Ȃ1zr��4���hAǉ�ӑ�Ef�6II�LYNQ���[Ե�0^��{<zс��)�ﭝ)'JM)-O2�oV�9]z���ɞ��Ze!݌s^�Ծ���2�k?2��Z/OE.tX��d�����dޗ�d+}wtAk�EpZ�#��[����.�E�3s�*�]!��0�F�j#�@w�6�%�o���I�7��|�>��b'���*��Z5m1TMx{@4�q�	>C��gXs|_�1_�f���({�u��l��1��P-�җ-�H������5�˵Q��� Ph�"\x�夣4@P�C<��Ŷ$gќ��)�^d�z �ųU�z�tY<~����ϱ������0���C�W��Nn�8tiȡg"�ecW{�|���Ң�h�z@��A�G�������K����1V.����:����ӱ���&��)�E3SL��	����)�>�rq^��Zܟ��o�j�#>�a�TA�Z-�C�K�	<��{��D�)@3�B
F�-J�^��p�.9�Tϭt�2��^�B�����]�;����+	�Н��7	����^G�'�y>U6$4�e� �S�UI��@��M�L
*�6A4H�$Y���B�5�<.΢%�ȍ��)�Z��{��R���������M�߻"�!��vR�۵�	ݲ�b�����S_e!}H�w����I�čy���YxpwW��}?�a3�>�<]�u��q�gkF���÷�G�z��w��~t+�����x�r��}#|6��gz�zP 0�U�Ʋ�D�{��t��?m?L�T܂InK�g�rğGy?P�:��i����.,�yē�S��Ȍ"�0�Ng�g-��j8>�UH�]��:�1�':5I6�JJ��d�ٽ���G��Q��$�\�¼��C�g�G�SJ�M�@��繌�b�<�SfH�Y���Ȱ�:�N����c��׀^�p�H�B-#v,X�v
IdRbw޺o����_LJ�k����O<q8���y�!�a��'�G�к�gv\�aa'�oc!� Pח�&���L
�Z�b�[3^i4ő�M�&�?î�`���>�ƕOy��!���տ�4�Y{s٦������6�\�wo�U������8t�p�N�"=n�K���|��z��I�%�
���3g��v=@54&Gv:ޢ��/�������b.\��#�q��P��a&��\EI3�Ӗps��|
N�	aT	h2��o	�-�ÜA��G�(��jH���dq>O����=�zM]g#��R2�W��?��ˬrd��ml�9֓ �!�=��͌ј�� �����M8����� �+Pϰe�i��'g^v�E�X��Na -��pu+��ߌ�F�L��f��9L"-7)�����G{��زe4�n%B�9Y-A�Ե3���r�e��
j.�}Q>��X�5F��rI={m��E�ע����!����(�f��2�����0j@(��&_�&���h֬�ժ�~1it�P-��{\�u�蝍YqM�p��7�#�MNh��Kbċ ���F��z\��C�8���=H��a����	CVk�{(�Moz �E���@������']"�)�X@F���#f���k�`��_%��8?Vc��W-*QY7e�QgLy���qX�g�Z���n\%~�"����ּ�c��^�z]ٍu�y�pE�M���M/�`���s�X��@��i<�c���^�Eq�n��I��9��5�?�R�7�M��c�P��߽p3S.+��|(�Wm�ǫ#^m�46qY�p�vA�U۟�������,��e�\YO���3�KFt�Ї��q����C�\�:1L��tקK� �2tdL�3���� ������ݬ�*vI��!�v��SR��-�PN�3t��3Q���tYl�>�Wɸ�Bƃa9�*�T�t��\�G1
�;�#"g��K'�����vb�#�w���
0��� �$�}�2��&�>7�}�$�
C#ѐ�ɒ8Q���@�p��e�Ŧ�)]w˾:/�[̦�p��-��T.43�(`�e�!e����96$1��w��^�gφ&��X��?�g�yy?��sT�K���G]߶��; f�u��+P�f���冞~��H��ukm��tՄasT����,�!&�%�0�g��Ɲ�8'C�fX�p��bhyt�)WJ�&~��nJ�]'[�ʔp=Pje�)-d��ȭ.�$+W��!t7˄�i��)�JO�^�͋�I�J��E9q���]����B۹�
�XV�7����a�=z/�49���:9S|��*�h�eH8�Gv�EϖUr�pa��^�#�;���e��ɻ�5W�-<
D��[lAsK(�������G�0���]��*ޖ��Q��l�,P����{z&����h�����(g&R=��5�{JH������N�#�x��2�8S���}�8mLZ2pB�t!JO0���F��ǁ��ߍ��!Vh&�A������Z�u�[�)�/�+��C�g�鷛�i[.-O\�YT.f�2���U!��ۺ��@,��D{b�cŪ�Z�A�6	��Ӛ�rץ�L�\6���N�4�վ����A����V���bBQ��&�Kh��ξi*�>d7�S�ޟ����9�o�0K��I; ��:�U�V�N?Ųh�o���b|9�ԫaBT*#��Ե��\k����R��/�Z]~�+�L�6y��'��(O��k�����d��B����D)��J]e���iu��z�Ģ��z_$n�K�
� %C
riMF��WTQDѸeA��,X�\r&K����-'p��T���u�w�.������q�����tPZ�����H�� P[_�N7����PV�?�\�>J<�-�H�����rHؐ������[zD��+�ha���َ�L�Y���j��U��Ә�8�%�)��t+ɭz��xy$�������گkщ�'B[��j4���c�����m݁��,�"��;ԦQD��7'�]s�:U��:�?^�g���CB����A(�F1����w��h�h��V|G��{����f'������=pu��~�Z{����O��~���_qCtd�'Xn鞧�B/�k���3�K}^Ѥ��t"L�c7�Y}�q��/c`�LE�pI�����ː5
ie�66"TY�n��sv܉P�8��d��0�o��ZH}Y�Ds�'����k,g�0�ἃ�V'J�:ո�����E�p�2���x�
��z��9�t��sg����yS�q���'�~in'_��z����[ђA�td�X9en��,_��i�` >�V�R��϶K��)=IN�2��O�a�F� �-���a���ݦ����9��w�o��ס,
���٫@��3�}���W�Ч��l%0ۣ`�k���Di.������;�U���Oͦb��WW�]DYa��Tqݍͼ-d��l���HGO�EkT����x`k�4v�Tl?˯�����v=�컏j+���¨N��dj*r՞N��K��U0�~�#�~_��m4 e�a�K@��(��6����S_x�PqZF/����b�����g�x��`�����+��7q��Ȟ�Κ�Ɖn��m��\���y��vM�����x��+ف�����0�ѿ� �r�K!م�;��q ����mBLL����PQϨƜ�ԝ[0��"a��䆯	r��Q�����P �nO�{�L`c��8�����L�,����d�Cڣ���B�mf0-���TPC��*q�����UU�ٴ]�k���YӇ�����`&7�����
��j�Vc��p�}4�W�YS��}-x����˿GBd��Ѝ���o���o&�_=���h�-*��M��JDY��W�M��{ZMK�\�-L,�ǣ�w����l�c1��PpUd�H�ڑ��~$r��>_�y��bN���'u>X ��|R��뗆�d6��m=����>�7��뿘�:�4]@�>���������$�z�<\IܽĽ�%��)#��X�%C@fU����sϚ���X��Y�g��@��G�^��rw6��s���yk �;�v`%��[�ߤ�S+Lٛ��f\�QbAlZ�;�:�B]����O�jp�V �ڕ׭�c��_�u�Mo�]��=�;�-0Yo,�����
�U�J����gI�xGxȝJ[��e��ݼA��b�t��8(��>H*��ns�϶�����v�G��1��.p�P��i;����,� #?�F�0��C��v����HֈE]�/�~�:du�
���x�����9�y�s`��0�x���O�����rɎ��b�{|�D��b�!��!��ć�Kf
���w���?;p(Ȝ��+�q�kӄ�A��j%�>)�^�+4X��C^-���"9���
r�S�+��S	G;0��|�Sln(nP=8���^/��PvyB �Ūʠ�@��c�' g�,s�����\�����+�TGn^0'~��XY�ع	�(3�ma�#��	�,#�|v�3�Lt*x-�:��}�İ�4�-θ�`W��Ԁٴ����N� ��r�(ۇD�meS�7��W2�7��̼nr��3�I��p��tî<,爞���=�i��M�A�>6	�Z:��Z+�1�S��a]���\�V�i�e\ݤ�����i�Cq�p�Zr����[��d��9C�����"1j�ʸ7rsU!F�78���%�"���b]k�,AC�ДwjD�~!��ͥ��7�(N4HO-/��j�*�~K	�������aZ�O�a)�Q39�cxn$�Hn�f�P!C�IaxYw���G���X?>��J�nm.�9�n��E�����.�R��=���Bu�k,�m�w<C�6�F����Tq��v;Pk�1=�h���{$8��[���V���� ��peO���(30y2�#��a�'��
�Ys9Q�;-�����7:{���L�G���8�n/�j2jzXNI_3޺�㜨�AqF
ٵ�	�`S}Nϥ�Z��?0�
�I9��͝�
��ӆ�С��@8�Hԃ�qjˡ/[$/��X���.)�����b�~R�Y3�$#�[����`C���Q_�J-��̤�޷�V�0a��A	g���6����f�L�Y6[;�^i_\�B!�$hn�\�J��Bt��'�4&��U�p����$,""ώЇ��=��_ȸ�J[D>h35���²� �6fOI�x%w�5��[J�����2N��K�Be����ή���QD>%am�i#{i��@|�`���ZI�q������2 �zl�_���,��*y^o�YE4�.8!R�o�ڧi!96����N�I�۶��Xl��/	й	�J,;�V�ʧ�s�нz �O��H8�p� D=h�%f5KdS���h�h4�9�J9j"�?�VT��u�A}��,�~N��f�f�P���
���)Le�.K{K�m,��Pn}����q��b� �����>�7�ݚ��JV��Jѳ�Qm�M��i���;(�i��帢K��7\��Q�1aITR&��x�$���R	m��	�=;ʠ���Y�ś�5�b75�Cdw�	O!�R�<����Ժ���k8k능����9_�뭌̴�gD�P�{��>�h-=b�<bS��I�1�g,�`�-(=h��0B�A.�J���kh�b�b��~�m-����V*w��߈M�O�~&a�\���ޢ����
Ks���;���0���2F]�Q#f4�q������H��9E;��F"�n�����F�iAoo��u66c�Pyrj�	�g[{��)m59��qØ�_;3�	����$����l�$<o,@#�o�9e^}Sm9������A1�A�7�}�ak":l,X��i��# ��E����r�񝽱���[����D�Z��;-��5��������E�?�D�:�?vk���2��M �6��j�����%������?��$����=���(xySe���[�����`���=�R�%�X(�`E����\dk���Z�%�1�gOHąq �LWph
�6#qR��ZF�z>�'�9q
R��I\�&?�KC�	/)	+B���5!�;+WW���)1����O��PaY�=��զ�Y�����T��?�o����{n�7��?�'I�r��2a{8,e l�7au��qw_h�?����'�HK����˞�њA��C�Oű7#	M�w���𣓶ŕ��R`�h�] �
ġ�@^� gnfo��LЇ�(���$�;~d�P�}�;R聹��0�u�jj���@�M��e,����z���!矇sBp調/�B�C}�fcs�D-����g���q|�X���D����r0`�q�x�����=R!\��dh�G3�g���|�A�у|��= J���wlT|�l�l��z]C���^��F��â��Ƈ<v@��a�M+�$	�g�W�#�4�X����-C�,6j����`�V��)������T��^����ږ�[»^��xe�uM|�f���ռfOs��'�s�f\+�?��@��_�,��9X(���HiU����Dmr�^p���b �Z�.5���;��7Ugˉ�@��&��BD�f��G���rm������F<���z�c�*��7M�Q����k�%{��Q�sq��k��5_�b�񠯥�˹�o�f���U�4�"#VA}+�	E=����mss���d_U��7�NE�"�1t�NAi�g����\�����Ϡ�oar|�D� 8JhخlR����s*�з]v�],�^@�rR���Q
4�+[D��\k�ʕ�g�h=���L63۶n��h.����i�͂�P���] ;1j�~E�4 J~ȧ���k\�Z�W5&��"��!?��C"�w��C%�V�~���̄���da��'��C�@�)�FrV ���n�)��iH�hs,H���WKܖ�rV�&��H����OC�Q�>z��2}|�'j���S�����U%�/�(4v}�Ҡ;J�x�⡮L���yf6'��A�f�@@E�3�iة�o'h�������c�bXi4�0��a��7���fEQ������]����:/�{���$O�C�YN��="õ���'�{U��K�j�SmJ_z9�a�E��|���O �F7�F��z������?�7������fx�om��q)�O����za�2ud\GF�����irzyP����\�TM�!��D�����ё������{���KC���\��AR$�����G5�U�,�r!O�$`�,><S7��~q�D g�>i�(���`�I�?1�f�9{x�Jis|�ۙ�V��#�ܦ+� �b8����cN���:G�&��L�!-)m��e�8�o�ܬ5�|�@4{W�]~��Z�a�X{�y�����3]�����c(��A�©�E����������!���M��G��g۴ǋ�h+t��+1AiY<pJ���/a�*�V��#-[�`�ҵ�����ս��]2���8��G�dVf�S��w���ǅQ���c�L���F�3�LN�Q�����=���@~)�պ"+��JF��IU+�5�+
�G��lԋ&�٨{�~ۉ������;o�&h�^���@n=�@o�Ib�����S9L�����c����mE;W�ɸ0�!��
T�g�9�9�-� �&نU�5ob���MW)�l� �+���T8vN�T��j���h6S�g�:�@��f��W� �}k�IͦTy#�9�: =(Lv�֒�gM�[�����G �(h_ >���N��@�q���j�q��l�w+�
�r����� �Œ���!}����S���R�;d��C栽�����n�����X�'�-�d$=�5T�n�ޝݷ�߈sB�3��D�IA�v���\�n�l��*�c/����^���L�Z��s;7�v�=��_��.ľ�eŕ?Òm=�6\J�w�Mbja����D\ ����7��.�K}-G�ު���9"�WB��+n�c䦮�{��������
7~�26'��oh�[��~�y�1��g�B�c��?���:T.dE���'e����tL�}[��;��6k����v��Д-Z7��F"C��� �����=��9
C��<Q� �o�� a�I*�*�kzz���*���Q���F���i�[�XY�v���`6�4�U�đE�z�Jy��#��i���;�����h�gPcs�	���-�c9���~s[J��.�Hό^h�4��3<�g5�ϥ>�}JeM��D
�^K���U�dmmU���M7,�GxhхMx��M����C�b�0�[��kd��#�+��tFi�~��d2� goa��I���8x�K�1]����*��
J�J4�k;YfQ]^2y9�d��xQR�9�4߃��\�xpY9ő22�M���rG��tу���þ1���0��x����%��5�v���P �8��n�����1k�_�b�Ũ��\P��v�V���\�zBm�(P�F�X���m��2<Q��Q�4`6n6��S>
�o�4�г�L|C3�3c��p!Cb��C3��i�%Y��L�*�&������P&wƺ-5w`u�-��|yT�+V�3��#�l�=�?:���`����L��z�ϟl�?�����ih���a��e��e�ӷi�#v��u�`L�p�S��ǜ�����O{�*8V�KS��"�~s`����- 2*�gn������V��s��@&�>�6FN��/l���2LM�����we��@#{s�]�FZyP6�O��$�f<�b�3MBo������~?��Џ�Ǧ�����'�=�0�f��c��^HIB��.^���0-�٠/ʭ����ŷ�3[?�y�~�؎�������F6��~^��x>��;<<���Q3�M�������Ġ*����X��]�/,S�x�"��NA1l�����B�M�A#VG�a�䪀��snk
|�"��7�@*U6
d�`Q���Hq���A��z�8ϸ�ݰ�Pi�~�McGF�$S�(!�y��y|	W���l��hdU��gBvuC�s��l8	'_�J5Y����v�8\�q �M��u�t��*�+�ǌ�s����<��K+������S0��8f���M���r:m�����Wi[㴧�3�jùX���A`&=QqM
� �}�Ì�����{�յ�s$A-Z۪�g��pF+t���"��:J8�`%�p1X~s�Z�2��{M��n��c��U��s����ʆ)�K;��"�\��b�q�]�ڽր����ᦄ��6����E4�q=�����=:Zѥ��ܽ+P�m��V�b���b�s�A�h�2z�pd[�so�'f�<���+LTj�ո���cQ�I�
w2< �/�+��0�]RH�Kl�@�6���Z���*���)�S]�Jo��8���6W�D����D���?X7J -��O$�9J�&7�u�����;��z$IR�Y�v�*6�2���q�{�<A|�S,�+R�I*!�Y�
z�7����S����a#��}Դ�ٻ���k�VA펝�~߈�p�[�r���6+�ɲ�3A7OMK�c� �������l�^��k8Ӝ�����?��1����Q� ���4���0�[k��0��o��[=�]PZ&8����fjỸ�vF�)������b�xW�,���[��ѫ���	>�k���.s�DI���]`�N�Ԡ�N>��Zr�w��A��;���T���Ű,Ii�s��ث`X��(����mUm�j03˲	���5x8�#�����G�4�F?������X�'2	m]���yLp�,rr�@K���lh����g�}�W�!�[wK�|��ʈ~$�-���:;YҤ��ن��	{O>��ǝ	j]�0t�Jݭ�knf6�~p���N�]��@l��z�WE;�a���yG�y]�	j��!����,��MޟL	Ս�4Z�j!���X�m
�B�0�9�:���?�P=�����R�K���\��k�L�WT�[-�}���~�@��_P}:�>F�vCٖ�9���$�7u��2�������'��j�ܖ��W��� �^�L
�HT ��`��.�%Mp��K���>Z@P�L�����f)�>z~?�jl���׊� tS��Z�t�����ʸ�SvZ|�v��HTl�q:N���6���m��W�hxgI�8A}�!���':�ە|h�g��n�kA���GzU�~l� Rˏ/������Ċ�sxz�2����J�w!�w~]	�꣸�o�!�l/5"��F�w0=�߸��"v��K+����@���G(G�C���Y�t\����`��-�V�v�F1�z��O|�%J<W�i䆭�8R�V�9>,r�J�&MTUL��L��҈۠}���N�⌺����)�4jKbSHQ*`�1�I�1j�g��A���p��Dg5 MċC� ���.huP�A�=���
�J�V��J�S'p�� k�=&�D�S#��u�ڞ���>/Z��Ë㌂+$���?]�8 ��֕ϕU{���Y��0�֑��%��a6��X�"/Xf�g����s���|K�Mׄ���0�%��~@U!�N*���7ofB�"����%�a��	X4���p�����i��x9��>���d���,>��C��!>��@n��lEY���$9QD2��v��B-����r�O�8���%$b���ʄ?X���,:J}3���.d9��23
�2��$XIwp�ly[ű[�>$��ܨjzN�����m�8�0��Z���'�K���j�m��{EJSb"��,h����Kyj�AZ�����^�L͋��kC�t�S�����{i�!���,C�� h�m�)�ڞZ\A���:�U�D��d��n(\��U���Ȋ�x�}��b�]��z��M�
r��Wr�;�͚���������"�ｶ%�-�0�I����X�l�~T˟