��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1�|�p�� �r�o�@���Ô����c̱��2�,fb�gGT�Fs�|�t���������-��xU�R!��d�qiĵE�}-g�	-�1���T
�@'d�5�����Yg��k�'���]�Ta!1�]��%� �C�;����#J\%mLܦ�X��$��@����n{��S���.�Z<�ٕe��pA�\���ڽ�"J�u\GQ���+��k�=�~n*�XE(�zv(���yi��?otzW:z�3ݼ��,7q뱷�����X��#QW�Ưi�U$�d�Bk�;�}���D0�$7�Z���K.�D��-�`���ߦ��9�7���# ��|n�#�*�t��$Z�H����I.��5&XNN�f	�P�1�?�]��a�8 1�1�u�[��u�Y����q{&��_vr#E'�NA_�-��;W��^Ow+�,��+ĶΦ�·!������z�a�yK,M轵��4cp+�`3l�Æ�~O���%eJ0j'�c�,�`�4���ؿ�[������Y�b�5���'Fq"������y�j�?μ���ق'�緜(8۰�(�IYxԞ_�B~me�������0��׻����M�)o�gA8���K��<�����G(���C�U�H�y���£ F�{���a�e���O�Yq*!�yj�Lf���{-+".?�h�����=H�쥎^��v�KP���jh���k�Hx��$
�Pâ,�ezU��I&H K�#z�M�`�^WQ5`�ܫ��)�|�W�k�I+�`ho�o2�쯵��,zwx���h�*��3�����3'9g��ۘÌm�U�8	a۠�@�Ǆ��.���-������%��:0$Sb�������I^���)�$	�Έ���YSɫ�qC;�b��R��_��PMCgxW(Is����-8Dk�Yܹ<�D�n�XY�����=@�!�A�V ���x]UD��3'���-�u\��,=���`��h*���a��*�*�d�(���'����a6s�&��V F-ɕ_��p��h��!D[�}������7���E�@e�VZL;��"��aUCu�{C���ac�L�$��^�����1X�G����c���Ƹ܆$B����Sa,²?E��\Q�̑) J�u���� A���1�1%�b]�����
���U�'��r>n�V��b��$9�d5����tY����I����y�D�W=vI�MqzI�d#�.{;�e<�*^9�ܝ�vf����>��e�̍	�L��F1�� 9Oh�ڬq̢$��猳0 M���?w�1��5����`a��i���A%J���Y�rU�=�U��`��-�d�1΢z𲢺3&ϝ#��4ۋ�K�7���PL4������� � �/�[�������~�\�<8����s�;�.B3��Χ.3�,7��6ug�u!�є���c��w9�����I���2�2U��+��xO�燈q���6��&@nM �p��A�cO/:�m�I�����ȴq#w��?j���#��saʰ=WI�������Os�P#�Z[��Ϩ��<��\�|���;nPM���m�(���@�4��&�4H���Ϸ���R�Y������<:�աSs��wdn�33�^�����Ɏ^����gǻ�%ӳ�����!��,���#R��"�@7�&K��)	��3�Z�ii���Qe�鎵��,88��|�2��Թ.�p���R�)jg�C$ұ��:�C�/gITS"BAQ�mQ�!����K��Ȅ����R�:k&�2�.[�Ҧ�Q����t�F��I� b5ޤ���'����*�j����p��D~A��ݑ'	) �y��4�<���<��%��ݿ�tU�u:�V�����������	Y�şa�ʏ2	��m6���"�u��ܧ�(��u��|/W�*~�*�6�':����i�E��X�<dѶ�Tu�bru-�O��~%���v>ݯ�.w�g���/6����55ܸ�y�@1�_;�1E0ٝU�TK,�۹	�s�������%!V�m��^���G~��)�K���҂RɌ��zt�'�{w�ұ���z 梹E��\~�L���ߓG2&/�^���d��ItN����g�.��s�/�6
H&�Q�Fq/������_��n'���igi����J@�kB�M/�����\��_X[������؇q��u�����eN@'��Â��V���k�Ζ�7���zפœt ��oc�@<�r�q���7��I��öֲ9nW���:5~���s����[��Q��˃B�G�rdPP.w���ab�h�I��s�b7F�N�?�%���(��[��V'/�6��d����?�B^���ǉ�S��{�=gգ�%���d�b��ß`X�4Aе=�rCF�S��ѻ������<'���F)DvpNY��3㦛�4f%!���>y�0T���'�!��o�#\�8��䙑,�L�=[!9ܫ��ffU���J��Tb�a� �fD�ݛ��P�┵�+�Æ�wDk��X�v��
ΉJ�ȟ����$S��6x�85������o�i�'K�Y��C�tI���ʋ���j��T��E8�a��~�7���'s�d3&o�MQ�����a�ׯ�>g8h�ʎ*a�Q=\z� ���srT�[�V֤6��V�@��X���I�񌅋�Y�-(SѨ����CU�m��
t�]r�|�E٨"͡��&��}8,9�1��T�������|\���OL� � yץ���m �&���|)PgH�x�u�+��ԅ* ��ab<��C�x�0��5$戀|p�����טV����R���,8��d�5�"^��V�a��*�k��d�#�aiQ:Ŗ3;d��S�a�{��,F#�AnZ�V|�_"���Rҙ�:_`�e,dZA}�'���T�|� `����+)_G�Ð�Of�/�� P�`y��^�����e@x4�NL�-�h�T��@xdP���P�1���B�O�����D���Xͫ3ߊ�!����L�k���	/p���_R�~�"G~�e���+l���(���s��r<�����F�����#��M����o7	(qnm�V�X�Mҽe�t?�i�c:�5�rz.�b�T����Uj��Ȩ�-ڟ�/��J0<���z��ǨP��x���ʈ>���g�Ѯ���z!��lp�W9�#�8���A?�"1��0��dd�_Yg�y[���\#9<���(��� +�W�U ?��vƧ��2�,�?fh�y{+�''�Ϣ<c���#*hI�/�O��ų`�明1�9B9p�S
V�1���6.�ղOF��6�t`�U�4�NQp�~��[Q�<0}ހoShy?�����KW�Eў?�������F�ŧ2z*J�Iu�7�	�k�C9�Zၯg5���UR��i���!|R���^6�]כ��!��\Z�8[��'�V@�n^���=|�쉏)��]�$����K}�������uky�"6^HL瞸[���9�2����k�X�]0�TQ�.Y!b{�e*�Hhs�\�MT��J�o�úZ�ӫ�r���NG�[_��q-O�E�o�~o�Z�(nCT��7�7��/