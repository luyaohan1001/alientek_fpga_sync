��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ����{��E�z!���o��>��j��_{*��u����H��WQ��8�z��-I�����M��U����M�u�XX�6~G�k��òǲ��0�<>�!H.$�3m��^�YFD3�]�������73���L��*���!�2�v�9Gт�"������-��R����af�{	8p�DD������!�Y�p�0	ed��SQ	ۗ*���a�v�d����~�S�65�LgiYE5���\E�{��9�稴����&l5�(���N\~��(�W�3����ݭ���I�X����a�7�H�����x����~��º�2�'�Z&��*׀ݛ�i�����?Dr�׃!Q��U�:q*3)Vsޛ�0)նݜ#?d-Sce�����3,��Z[D0z�癣(_�S� �F��9@�h��B��b��X��Z�"����R�X��8|Du-e�����f8�����I���r��2;v$������NY7�A5,������,+$�K%T["	6��ڴ.#ƨvm�����ߩ��e��dD����Kx�!��~ơ��L8HJ�V�rq���i��=z\������Oҡ"�*�Y����r}���*K^�}i�N�z�"$G6��Y��t?�Ŧ#Z�C֒A��X��-��q�K�t��7�2���p1QL����|i>G�/����#]���s��/x�É̉|���+�0s�2��Mk�o�U8���7�d�lj���<1Q=H�o`&f�5
/.�b�1�^�˩gF�J.�*���t��.�� �&7��S���h��ܣbD�J<���W&1 ��:A֤���.�3��tt������G�r�JO�����kx��u²Xv������	��2��Sk���0bw�l����m�xN)^�i_���c���&�������a��u{�0��A�%���0ۼ7JT��}��l�x�^ΐ8z��+_i�����j�3p(OM#F��x�:�Gr`S���x���KY7W����4^Rc�#�����Q��� ��]�n�пr��+�P�.��O�w�pꠕ��T��T̽|o��ؐ��z>0L����0��� ɛSy��j!�I���-Q��#�hC��E���lđ���ja����Ix�i�jb�K]�a�C�ț����yWNP�'�����Q���抦ۏ�a}�X�k�r�n��Q����^�1^��_9,ҏ�E������*b������`�< �ߚd:�'��Q/����%w�"�f�
YR�$�3ړ�"�4RLwl�q�x*L҆Q�T�S9R�%Oҽ'7F�`�e�R+L7�y��"���R��0}��[k-C������0�d�J�iRiGᱽ��O.'�L���0�S�4_���Ą��7Dr���|����@�9�M�+��N�*hi�@aUC��g�-�������:�Ch�rm뙮Kw=��<$>�
��CE	C+q�B8�x4������Sޘ�Q�u��?IW�\4�G�Q��u��� Aӏ�$"�l�V�v��z�qR�v������������'��`E�oB�AWǌe7�턮���h�N�r
?�s���{�FU�q#��`� Y�2�ˈ:��������� �h\�WtVT:#҃|��spإS��*�֣�����Ah�e��w�2m.ַ�9�����4�;�Կr8�ld��c�Z`�SLTc0l)ű �	��~SR6��w�W7O�I��8Ir����g]���p�N{����;���}5Y�]IQ~ ��<�-фk!8�<��p���ǚ��P���#��F�� CS��$����m-3U܄����w@l9��@Pw+�� �c�|�"Ʊ'$R��^w`_�*�z"��Lqt�_��2j��(��oW�!�q��rC�vo�;)΁G�N>_�"�3�G�#���B��"��]�te���k��48�M�	a�V�:��9�߫���Y��X)@?G\�?T�ӽQa�c���8,�N�j����E���R�n�;�[��,^�n0��v]+������@ko�6i�82���E"V�!�<u;�Q���=aWE��iު\!!b̀��'�h�@����� ��>^vp7)3���6͡U 	X�m�����g��x�R��	���(6��?����	h����(�8���3`�t��!B�	$��ؚ3��O�R�tQ��C�f7Ҭ̰�^s�w�;�`���1�2C�TyR�ٔR'Y� ��į(�4_�7r(<�(���Fm�j�������b��l7?vEؖ�%�ꔈ��S�ꪊ�
U��G�3���T��~g�	া�o��'|����])�"�W�F�-j#�W�m_X|�!�#�f[��8C��z�u%����T6�j..�r��m ��Җ���]��a�b����[v�SO��>��*�a�O�4Wg�.��^��"om%���?����50�����:$��7^�(,��x�	
Ni[� u�=����4� ���l']���" �o�ݦ�.
T=E�����mXXY>�؇g՝A�wz�p���(����(Y�[%�׮!{@��:v�O O��	�zMz�%�*&��M��Q��L�2w�Hc{0@kH����5��Ǝ&۪��S
�PV�����4��f�s���l�fֺ�BB,.Ř#����y5N���'`(� ׫�wX�)����?�㺽Z�#{�Qڱ�(<����?\�����eI�����D?��Tܧ\��C4�9 �	�q%,O�#��:i�B�]ýZ��M�8( �O�{U�D��ʧ��F�>n���5o�嬤�#��ZȆ��:02 BE����ә�`��jX,66�L�q�so��r���S�Ǻ��c0Tp����Σ/�hƷ�l1s�W ]D_�|aKT��� �Y�h��o
�r�^��Ca�!i�%-��M�8_����&藼����O���,<%|�<�#������ΈIz���%O����Ck�U�{SGr���K�\A|��{�z�]�)�� ��"&R��>�>N�^��r���&�Q��{$�O7����3���!#�%���)�	·
)	�"}-y��	yC�ߴ�Ғ�-�*-���/�����MR��tB�:�*���MI�>�(�&�Pܗ�L���x�?,ѫj!�m	��	����9Y$9��x�7���p0n���U;��G��#�3A�٠�n??qUK���oY���]�������c ��òq�}�]���IS`���� 1��M��s���x�>������Մe6!��\��"��&�Lͽ�� Y��P�S�y��Ϛմe���b�d?DB�s�2D��h�Ժ���������,�&^N�����#�Z�m���z3Fh5�xw��-8*,&��E
��+ĭ�
���y�pR���'Q���9
���3�2R��k]�i��K����xz��P����v0�9�(�CF�¡ȫ'ә�ڤXF}zĺ�W/�5�9����jJ�~|ڙ��"#�C;�$ܱ�;����b���;��zE�2Y�Z�m���3_�Kkm�&¬}g�P�p�p; MvF���;��m~ݠ���ȃ�6�g��s<�lg���1�%�2�f^�R�,{�/y�:Tb�G��a�}����򻽞'@�K�e,j
I����2Rrw��H������D��ts�]G����+b���U������ٻ	���=!T�^\n���GDɹ�_���R�I�?�I��2��'���+Yk�!�p��k>�s�w��8C��~V'�^d����駖�X���N ҆�LěI���	�C�b��[&t��f�	��m�����)����e/��v�Fl�D��>�tWd{��`��<3il�y��?2/��{%��D�ȴW�y�n5Bݺ"���q�-)��g��7�A1()�j���ކ��m;e�^��0��n~l��s���u7�q#�l������v4�S��6q�Գ	�#�FI=�ꕓ#NÕ�O7=�/�8�]0��EJ�	�z�!j����H�R���^.y����3�V�I7���Z��6�XK���Vi��iJ����)���$���"����r���%*C���eC
n�=��I^(f*��D�4��y{�D{-o��M�<��\N�R��°k��\�>��}��&�v���!k#�?��	�驷>���Ž��E����@���S�?<s4��\V��u�T�qK:s�:^�#�L����f Jy�����U�,���e���S<�m�Z�"8���Wz<��"����m��L�OV՝��'ou#��5�k����2��%(Y�&p�kV�F�˅"����$A��qg�߫�EZ�%�f�x�DgoB��uQwF�0\���6�Q,�5	-�6&�ʥ����
i���Z)�ϛ��m���eA�Df�U"Ӈ���&OQ��b�r.��( �ą�:��y�Z>p�NOW�,��8��W��3"��H��K3�ϡj_D�8�A�j�_�2�@<�@��A�yӑ���L6�h'Y�`|��t����M{�Z]TA6G3L �]"����Iъ�i����k����F�2f1��^�۩68����%b�q<s�r�el^@�����ߊ��}��\5T�A�;�0ѼSs5B �5G^�����!��M�����H@�hlH���I������&����eEǰ-�W����#���g��
߷Z�ҧ����a���.�Sa��f����<&�B���ƞd��d~�wa�D9Ϋ��5f1Ec63J����n���lD�Ӂ �9Q%��n���;u�dxJ�dm���oYl}?����L�����f�0�O>��^E�x�I�O�8Q?�CU7�6$�JH����ᐁK�ѕ,���Щc���![:S�q�i1���"v��Fa�<S�'��T_�_�s7��;5R)��2q�zd�Q�z�I<n%o|�Jw�[��·:l�W����S>r9�r{}{� g~�t+K�i�a�~���m�9�Bu�vu����n]�r�;!�xO����ϋ�;���*O�
�"*���nZ���[H�1�%����̊_ͪ��#��?/�nģ�a�m���Ҫ�*���s�ik7�:�]��z\]k�����M�E���<ˀ_l[�2P,�T8����7�#��o�|	��V�4�2%W��āu�2����'�:/֘�W�D	�6޾bh���N��C���֋�b	�K7��?���V�i�t?�1���h����D.1=�Q`'Ū�"C�H̰F��!����d[T?k'(4b��=�<�}������u�Ѯ�Cؗ8ͼ�����RBZorL�z���:�h4rGBR�w*8�V��'� ����~��l�Pa�=��^�x�bv����T�v��j ��ճ��|�~R���$�e�T�w�2�����N���g�ܥ!�ú�O]�4�B�`烙K]Ѿ�ٛ�F��ͽ���� �qX2�"}n��S�]�� ��+;��������|�J�㺀G0���نs�P�l�y���:7UHP�a�y�F�!X4�	[�J\��ý�L#VOXJ�=���)#��d��H�C-1LK��mkզ�;S�G^����Yd��Tį��{���^Q�%�w�%�f8���3�*p���w�!fq��E�_=�$ ��'�6b|"���_	
�lN��<bv5�� (��K��<=F�~f�333�F���\Wm'F���У��5��<����%EA<���~f<7����SMRZ~�զ�ߧ2�Ί%R;��`HZ�Ԫ���@g�{���o�fU7?	��Xh)�R�_f����BE�D?}p����|ÉS;Qa!:�(e�5����ѯ�oa
������HA1X �����%� c�� A:ab�,E�&Q�d�|��5��V*��˄�L����@f�
Ha���Z_s�c�{�Y�L���ܟ�l��b���v�����Dw
�n~���4I�܄������GĴ���u+� <�c��XYQ7˿�8����%e+�\҈4h��� u�Q�g�ӆ{ }�N�¨{�`0e�.���GP-*&+�U;��j�(�A��36�yi�w�r��Kt�.�~�H�Y<�H��I�y�<|�ZcU镌`�m-�l�>Սs�洮:�)�-D�7,_z���z"���	d�ߞ��M�|(�6s��yfh6�Euʒ7�ӻ�����œ�kx
dr �I����)01@�&a�=2tP2��6��;V����L��@����@��e�G�����K�fۥy������p���0A��GR����c�F�M���UF�7.W�s@؞ি�x��"�$�8|��aO���+�`{Rㆭ�X*���@^��,����ˆ��`���:o�1��~��
�>���J28��)�T$�q�ؒ�mn��hYc3��_��K`��J}�S�G'�M�~$���O�{�nw<�q_�>ٺ�|�=*���%��ǋ��U3�s�Tj����C��h�D��_�d
����68�CG� �|��<b�����E���y�0&Q���.���S�ţZC��p7h�3��Q&8�1+��8>YE+R�����tBa�5ȼq﮼y]���L�;3���ޒ{4�w<��b-��+>���z~�T�D|{4����2�C�s�V3Ht���TN��:6��N� � �b_������O/�Z���N��t�ls�"NA$����$N�2��ee�LH�\*�Jp�o����"wd���q�Y4��~��c��;?���Ld�X�?�?���eڗA�-Ip<�=���p�6��G�g,|7��f�x���Pm2�Ymkm/Z4Š��v6�|���0���\�l[y�ae)%���a�x�4=�����l�_x�4A=o�qe>d�Aw1���F�n�P��Ñ�1Ѕ��N%��5�d
�1i�ċ�Y�"M�� 8��R�Y�A��t*�.
���I/N��n���\�"�0 s���)m�/�m��&�_o�K&<A�Ac��R.ܚR�I�)��b���5�e�:׃!�
�R�����_�����*&�etM'=�՘L*�_<P-�:U��A�!�jg^�^�}T����iH������W2;��>.���wE����$��]���c��Pڊ�4�z̓���6��h���}�A#{��S�|���E=�l+[�Qx<��$,��J� N�p�҃��*1�h��Z[�џ0s�,m���x2�nf�Y[�wB���;�_ڮ2�&ޯ�NE�>;�+��S�U�I�����?z/v�V©1B1-s���$"��h3��߽�DT��j�p�Ji�E�N�����}���B�7�.�Ū_��
Ƕh��mW���B�	>��H?m��
?a5!����a��`RP�kP�ޚ�H3�>��+��q)��GmG�J�+st�I��@q�ّ�-{��n3'x�j�j�h�G]���H�Q@k�_WX��ZbU��8�RD/]�[�Ti�`i\�-�M!Y���ta}�ݨ�A�&�E���'�Q+G�k����\�іv��t�'�k?��K���EJHO؆���l�,P��Ui�k��0�!�)�x_�W푙(�������q�����:ě��H��(3�W��5���� R��G�2͟AM��:˼g���cEǋ8�k�,���m�v~֪���sc�a���c�Nћ6���F9��vƽ#��F%� �lM���g
�״��o�U�����O��Ļ���1����/�I�ݩ���{_�P
9��v����g�`<?��o��=7��J��J̍�{��{ʉ�"���A\��.�Y7f�����.�Ϝ�a�q4��|3 E���}�!�9<�p�_ U�I/h�n�8��~�trfmL74��h*��B����yM�c4�A>�`��޺�ݘ�}4�y�����V,f���-��&��*��\�..V�R�8���Ɍ(�S=��y�ҘTb����d涡Q-Uhʫ#Sz�Ư%�=�=�FN ��a�#��Էa;n[�v��L��a�n��Y�+��$�?�L�4�u��$�v�U����3Gm��a�~��;d���F�q�:UI��x��ݎO�;��m��\��)��@�+�]Z�ӱ������cK!^ȸ�@x�TşfAJ����3��7�����U�Ed��d��"n�Ruݕ�CzJ��W�.?���FT���f�V��Lu��9��>2|ȹ^�fUi�
��oK�F>��;\3K�"a��z���)Ǒ!�E;���Ug�J��.m��I�NĖ�xLϔ�w�ZVh�oF�`� ���M~b�y8RYU��,6��?t��ף�0M����5�_���'H�'�Zw�{}���7���F'�]񟢞�My�x�^m H��������q��V��,�M,+vָ�㕮>�k)��C}8��H�B�{�67m�v�Ԋ�	��)�C�6���:��a0��C�<?��=۪5��ʜ���oU�����o��4q��$ʷNu��E�~�lĺ˺Ի�c7�ǹA���FS���G��I��M��jw�{"�0��v��U�Nv��P�ܓa���b��w�G��̨�l� p�P�4J7ye��洀��]Σe>:Z���W�	�d�U��p�"�IR�;|��s��t��ġN�����>�&г��ƹg���J�}��z��	�3CZU�5Ͷ4/�!vYB&:�e����WyN��seD��}�/F�;�b�c?��gl�d���uJ�YR�w��(Ŀ�K�,����-u;A��e��[g�^,>��?���_��*>J�Vp�
��x��]-���ne�����Gҷ�Ig0%���X��^'حv�[.gXB��a���lg�$b�Z-�l�@��rV���)�^~G%}n�r���D�_�P��xu�[c�y��{e�z�X��A�|�����[�9$�.$S�~��wWP��Q�<� �c���b����=h�Ҭ!a�n|K�q��'怟R�Wr[�ev�0+��¼"}��x!��o�FT��V�DKZ�Pc���AK=��rtU��kr�c�m�O/�#�*�wM�&����QBv~n'm�Cܕ��/���+ө����3l�� �*n��A��A�z�njJwƞ�����#���_ܓ�����g�g��x8�3��OUa���%�˛�ѠdW�E��N��K��Onv���4��c��N�1�;�uЮ�]�O�!�Ƅ��碝 Zm�Dj�E:��q�8C�I�ed5ym�9יQ���>�,�?*�w4��p��XBe$0��i�}9�n1��C���&����ϡ���Va�5���+q��S$\Q!@RPe�*��+L�LtE�r��uHd����c�<�r�>�f&������C�p�� v�A���Z��c�'��.N��-12�2АE/����R;��1��M7�C�������*m�N�Jxv�l�H��EYC>a��j,�� �M��"����}��Sl�`���J��M�f5�Hb
����ɝ%zѰG��`Hk�/��k{oqs���������G���My5�W���	�W�sR-`��3�w�/��y�h�_�O��D�z�s���i���mE�/���ϕ�bV�I�b�r1��?�39ɑ�N��:��wu82� -�8zo&�+	�o���gj�]�@��p��L�0{�2���6Bm�n�Կ�ٚk� &�1�cUus���v64 ǤNF�y��+���Ư>�h{�S�E�Ro7��+ٹ��y_��*T. L�
���_I=�јK=æ&5Z��x�K0��X���ɱX���Śq�ϒۃ�g��ac������Ȧ�
�����N��H)b�|9�₏�1`�vi��t_m�`9�N��$�2�^�I������Uu����h��=�I�3�m����Z4~�֚�=�I��x<�p�V�/P>�d|2݆!���D����{-�p���%(����q/!�Ⱥ�W�8�⏋�6�'!�^���}���Pip�-E6@��{�6���	Qv! �-f��O�8^�C{�E5�s���C��*�Z���Z9T�������i�Yc�@���S�,��m�=�4�˥�7T���f$���%���ѷ�M]j�4L�u�K�R�YG+3#0׻�/�-`���)���xTґyљ��'���v���y������z���z�"o�9�
�6�@��wn��Dܭ�[:@K�(��{ZZ8�.5�qK���=���}���7�p����@���J�~���B�`H�1��5�>�7���%���$Y��eח�2�E��u��t�0L�{^G����f�'��@�7�c�.�������j�g�0(���a�ïbe���U:�.pn�G�ZrN�n��*%��?Ta�ez�e)�4Y��Nڙs*_lݿj�����b�1�~����yD���`�..l�Wu3�_�B�"$��C3ߨL���/��P����'�n]��"��s�5����1�߄��hݼ���8���Sظ�hp��O�f���ՎG>MNGfl	�9�3�������([�����!��EtX�Iw�F��;M?[@�R��?���a����vg�Ew%��t|���M��i囘f$e�$��1��F���M�8P4��>�.�8��j#uō2����3��ގ?mR�^=�^x��=zd}�[<H�^����@�#9�q��7�mC��`��%�m�0�Vȧ�:��5�}�y#���pVڝ(����o�a�j�S��0gH3�@�т.N��I$��Ę88�a���E��	t�h� i:W7'[\ކ�$#�OԀoLf��ocǜ�.:&ĳH��0�ݡ�T�����/`x�;`l�����07gs�'P`Y7'׋[p�@2�VK�ן�h��������oU�:B��T�L61��j�N�"�9��Ul�b��r��=ڤŋ8n1��y�Dt�t\����p͉˖��@�X�E�[�(��H)A��x�B��ƿ��Jsenp%�%u4`�n:�m��]��3�2`�\��wj���q k���a���ՁfP꼛LĂG��x���q}L>�����5�
O���΁\$��0$�;�1�9օ� v���2�c���!�$�!�"%#"��m�9Ͳ�h���=��Б��^d�W�mNc�>��8�P��t0I�3������e�c�?�����=ť>��
R�����Z;�`�{���a8��5�d����{���U%��e��T�o�H���P�.+�]�f�� ��Q؜ �;�rZj�=<�p��]u�7�s~���3� е��	l53`�)��4�����$Z���_�q�>�s�V�\�a��ma)yM�@Zxߤ�|O?�����@	ny{5Pw�_I�6P�)�T�x�X�<�7i�'��*W�+$,T�u���R�� Q#���;�j�@��)J C�{E��t�,D�ɠ���Y�UG�3 n.�Ǿ�=r�<󯹱��4%��T(���jf)b�l���Sy�C8ʨ����a��x��t��hh)~���l�"�/Nt${-a/4�lN7��}�����<�1�[ठ?>��W	8=�e�0DNΥ� C۾d��%��GR�Z�}S��L<	�������w��f�XI��b�����s�Έ�(VmUÇ�Ֆ3�t,&���GYZ!.�����"-�6� �Y����p-�m�~x�S=�����xE4,B5�G�Dn��I�<��dԋ�y���yK��U��8Q0LL��2i�,��|�3k$�u�)>��r�Ge�(�KP�r�<#g��E�#?���\җ��9�V�MU ���;���M:C�Q$�ƻÈ��B]��7�K�#<�w⑗�~,s�/�i��E��̮�����]�k�s��qr�p�\&d�E�p�ެ���#΃���m�{����tXh�/<�%D,���Я_?q�޺��Z�������%t2��z?<�U�]@�5����O�U�qtV�mw�&bن�����n((�榴7��
��	����s-f[�z�䍁�Z����@���T�m1��~6k�p�{�V�bU�:���)��@��X��NM�Gإn��6�U ș�>e���#y�"2�%YE"�~���9��=y�I���Q�
@���a'	֗L�
���ue1y�.E����J{�<�)�� Y���2�h5�1��զ;�|W� Y�!�Hr'D��S�¢(
U� �h��M�V��oۙ'g��I�`������ �S��7�axڳ��|���J2�9l4��/���ݢ�w�b/'̛�s=��d�Q�r��VK�?/�����pS#\��6hhW<a�h|��dyr\Uh���o���'����3�J�i&%���5�w��4ѮyY�0��6�������QR�z7���!��G��&Ϝ��lNJR	O�,� �1����2k���9�,��L>�[�+wD���9��C�����֩�y/q�z;O�X� CD��7�頟�K.�4�	�N�G,�n먏\�wB�i�̟�nI��������vgkkXu5b ���U��W0P���wQ��n�V�U���ω1�#뤽/��\{6��~M�p����,y�x�o���s�I�t�_�]MX��������tP%��nG��2���W#�]͗7B_�X�G�mTI[���	8��;X;�0L]B�k��P�K�f�o�@���џ��d5��1GWs��vd>���O�Q.�EWJ����K��#Dv� ���S0~F.z������W5�Ϭ�vx����|_"ە~<�?�Q�Q9�_�����
�;r둙�)XJM���Ғ�/���̏�4�6���-����r�TT�������G��	g%[Mi��"�������n�)'���O�0�s�y�	�U7_��$(@�@H����UB9�)�I�� *~ii!����Q�Bt$$�ޥ�z��X1���F�\ 1$���1����(����
gF���+o�j#��aE	z�^d�tC�v�xz��X>��i��^��n
{�������5��K~v�OE���l]�	x^;ʓ������m�N�ິL�c�aB�2�_��{�@'��;O��o�?q��P���\ٞ��\�<����+\e���ƴvY�4��S�Oߎ��O4C���{�[��R8���z�z>�F�lF��4܉����j�o�޴�N	Q�ds��')bdMћ���P㹼ѹE$>��G�,�\D�j�
LT���7���\h����LE�r��ש� �_���z(H~�"\��]�;b q0�{@�Đ���p[�qM�զ5��<|-�`�
�W ��N��ҽ=H�)�¾ˠ&�}!�i��Ǻcx���o���WSi'�.Q�j?�T�s���"���JM���DN�����J2v�b�^��B��^X��8r8^�ǝ�,��X4�\A)֩G���н�P}y>����wb����w�b`�d$��E��Ip��Pi���� 2 ��h $T�`_/�(,\�R-�zY[sA�*4���!8���@[��:�5�-h
��� �>g�Ҫ�Z�f���\-�>��lv����~`�e��u��9�U�
�pp�Z9A�(��ӳ�y�I�>�N��m���(G!Y����I Lʭ(8t���M�I���y�c��&�	_CO��b�Lj��r`Q�N�^�&pg�i�	j�	������M��\���Ch4Y�Y�����S���}L�ݲcL�=.Q����xz�� �=��H�������*��>�K_���N��E�[�	
��Ф�)9P&�+;���:�	Y�G�]c�z)i��|���먛����]s�e�V�`���u��@Rf�iW�����W2Dww��δ�ʎ�1V�v�U���s�������	}�|ѻz�	�����t5�b�3*�\�����<k��u>��-CH��S��A���od�߿!��,A/u��@!\� y��9�&��a��1w?t���a]��?,�%a<�|���5'��k�FgV���Hq�5(b�!��4P�0h�*�G$.�n`�(;�\
W��~j�r� 4W����C� �-��u����g6�J�@�X�#}�(օ��hJ��W�H�հ}I,��)�{�<*?����G�&͗�[F��(e,�7/�"�����m��nc���Lp�g�1����g�{�[�����z�ͨ1�@3E0R����*�}��|u��#�R�,afy�4�tK����L���Q����V�8p���*�i�2	�E�˯����])�n"��Ur��ffl�$:�o� �#j ��]R�H��_p����	5&���wm�Ύ�L����W��
v"��7}��2�v>����� �o�Ơ�z�A2�5��� ����aה�G}L]�0��P��U� sⶸ�_,%BZX�(�0we���/�Ea���ɒЕ���0�U/��8�g���6�ӷ>��V����|��r�g����\"�&0����J���Mw<��O���*�����5��:a��}���i=f����1�����V���0���G��5ٗIk;X-=���P�mO����8L�MAtOe|���
q��ۈ"�W�j��HwĔ	�Rj0��B�I�7�!�%�R�$"�/oV5v@=&���|��l9ˋn��e�ں�k�`��uz9�9��[���m��F�]��:'�Z�X`�E��U?R��"I:.8�G<�$��(�U�1O�7l���Rk�EPnPY@��՘�r�p��!�!7��⾪C���� �gp�bG�YM�����:K���+���\�2��z`�
�pD�+4��E�$�b�Dye��A7�Cܫ�E�q��m�u� |��7^x_p&m�W�=��3CnJ�/}F��2-Lx��[�r�d���a( ��TOő�P��ǣ��Ǒ�b��O_�ȅvL*�rᲸy�u�-z�K��Y&�w�����>����k� ~�@��� B�4HB�	�_��g� ]c�BF+R���Y:)���LI�[]p&2��2=y������Z�/�g	֔m��e�MmҔ��`i�1����/S�����[ʈy��}�}E�b?�|aZ�����Q�X^ڞJN�%K��F��}~z�^j̀�<�T�+�]�:�$������~v�+U�籌��{l��!�d�8K_ܞ�"�7�@өT��Ѽ�Ξ�N+���c�.�o�B�L�ހ��N-$�Tp��r'�(	�7$Z�r/$�ҧ����-���,�ei�(��Rc������\���2	�_c��eh�/���e]"T0&�[5ڝ	�ma�O��HI�l0.˩�c�g��x�ud�Ҍ�a�FϜ�?5���q ���%ҹʼ���-���C%��J*�J���:*´:!��_�\�`h������y���o眩ҿZ�/+�L[���m��l�2rt���;j�g�Ƞ�[�P��������~�no8��#&7�\��S�Ѥ��?7�[��"�{�4�V��6Ͼ�>H���7��-�~�,~U�k9Th��J'Z�?�h�2So�U���ȞH��?����鯥V�iG/e�2�`I����������D3U��-zݔA����]�����}!u�U=���U�/c���Q���pJ�\����l�/TC����G������0����S0���9�o��Y@�x�i|�H�E-�GW�Թe��h�;�{}'�#Qz8���u�aj{����iic �"�ORu��� )B1+t�T��n&0zG��7>���z����a��K�0S ���+u6�����$ p���T3�����^Pq���r���q�5d�_wc�O�m�{ܓ��&&�ǌ\����S�_��L:�o�0k��ͮɜ}�]��y,��z��������t"=˲
A�G�8���8*MC��[�ީ@R�n�o�(�g\n���������H���%�;|:��c�ܬ�~&s��W�>$z���tg�X_f�=l�}�9��iL\m�<��-�H�R�P��V�ޡq��Ӓ�����=�6_�Ux�� �,_��f����%'���A!�k�E�z\���%T�
��H+-���̎Y�v}]h��K�Y
��&ӛC�0C[�*az���bR� �++��d�h��z�)���i����N��o'w��<*g�^��9P:�l9;�i�R_��-�
���QG�|B<��oW��w� l�?��`�дMKX�E��=@�ƌ�~4���$�.��B�=|;�_N��N��X�4>��LZ�?*^ta�j�_���&� 8V��d.`>j%��I���*��DK��E�lH>��h��~Q���7x� n�\Bќ����4e��5�� �a��9	�n���/pL?��jN�$�+S?����fE�a$��S{Q	�"/s��\I��]��}��DF�m�q�F ���j̼�{?B���^�!%��K�(�D����tU�9M78oi0H���b�{��c�|�����;�*_B�u˿������z�]�����]l�b��7�-r�`�.6H+��*_�\