��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G���'$�ƣ�@a�=p*G���z�Y�%L�YJ�V��t�(�]+��ZiO@��l�2,A{���gA���msl�T�D^y"�h`=[k��G�4�/�)~��|��O|�5�9�����ǳߤK�韝��	z ��A��7}�+\�`�d)�F"u��λ�5��u	�y��cy����|���n���h���ص|�]�%ߨl����������Z��C/�_��P3mi�9�g)���i�t����$,�d{�J�2��3c��Z`���v�ī&`#1���4<���kK�\�)�_�ZN �'/��E���c7l�3�gHq.JK��5�0֔�Su��m�{����}�9�|���h���[�H�'�ɺ�r˄��_����W�:�\��Q��o%jk!�		����@'�u{�K`���dc�ci�٧=q�s���jo���3J�Y�8fk�d09#�8���y3q7茹�J�*V���M�{�gːA�T��M�Y�A������$�IO��SlK�.pR�|k?��6)bM�����n�>T�k�{Q��C��(�����W%��pin��͎���"��=��ȯ���#Чr�%CvBS�s���P���ϭ���TE��t$3����Nu�w��	X�[Xִ�u�n	�MY���W�:��ӹ�W�ظx���j2��X�͂��b�؅��$A��_�@�GA�Ҵ�ܓ���=�$M5����^�!Z���/��Zc��_�$w���j0����*|j8T �����n��V���	�k�T9��~$�����)r#/��ȗ	o_��lo<��)�*�aH�؈���%�]�S���l��^ �����c�.���H��F�S:��"��ɧ�t�g��H��c1��v�'�Z�$M�a���`Nf�E����LR̮��B�q})�A�X�{���k�P �N���U��Z��@�&e�<޵]����K����/L�2��}��F��s��i�����JsS�!�K)��ː��s��4Q�׳�S��z&���ƙ
����qA�A$|L�� �̰
�`����!�{vA��撌����^�q-���^�l�P�����	���-�XR�·x���̍Q/2�c�,0Շ��"�Ug��28�������O=1�0�%���-hCxaG�,ԪO�w�8bQ�W
t �I�gx��������Z��)����r���%.4��~�ϭ�¿�h�E)F6%F�8c�,U]0��D�n;�n�>y#�:��	[F!_ggK���n�m������mI�O� ����Y��&3?�U*�U�ڣX�g_�@&�s	�~��W��(�>b�P�XV�]�7X��s�@}�I��op�A��r���b���출��:�[������D'g���H������M�Y	�\�S��0R������0E9&��¿�o�}7u�HL�ypH��c�I�/��sb�\���_�ܹ9,kj�kG![����bP4�����������h�b����#+�/�P:�KKc^c0�P�58G.��?���q^�DKT0N1�(N�͢�ř��)E��NoO֮�~�͓�b��I�] ҒC��K�m��V�����XT�F[��3!��	�85��X��^q���m��7tGn�oCZo�����%ᝇ*I#u��3���m���&*�i��ۺ��_I:���~���\� Z�j�i���ZC�t ��47Vz�m�m��}	�<j:5�!y�7��)3L�ߛ$A��بv86���������t��s�P�t�U� ��`r�Nv��o��v�̱��@��ճ�wQ?��=[G�ķ��`�`����PD2Q��_����N߳8��%�&�&c�v��ژ�!���xbh%�'ڠ�aO�B��XrE�]C�}�9���%���b��EE&�&	w�e�����:�k�2u(���N~��2��K��~F�hi�˄X���j883����R��,�b׻�w. l`r��i��YH�0WsSy�E�!Oξ*��=�O$��ϩh�3��߾GF8���f�:{,&6���"�MH�oej�V"�	<���81���s�ŧeO��O������@�*�tS[F�1Yv*ZB5�v�S}�L�.��D*�m�� 1�����W�����o��߫n
0Gp��_��6�>q>*;K�~ܰ�0$�(�1�8���x2J<��%���Z]�*�,�V�]ʣP��B��zGX��� u�\�Z���dܫ�`brԅw+`�?I#�Y}$�R�(����oD=s����c����C��Z�I���Wr�@��F���p	z�o����,�	�̚������rI����O���Z���e�́�*�U��	ٓ��P���=x����콅Ҋ���?;��_�S{D/�ҧ�?�G�Y-'��(z���y�0	���G��ҫ���u
��vXp~��n��.~̛
B^Q�U^]z�.�$؆}�y����)�=�8o!r�L?��W�X3�>��n��p�.�@B�cΈ�; $MC
��j��9�����B�,��{�jIU�]���)<@e��$^��Yl�����|���_A�F�aV�#��
����M}�o�X��[s�n���b5�8�6'J<<șv�{�Qb7�3��^P���4�m��M�|�)��mLKm�+w��R͵GJ�=q�H��aByȕ�8sL�"tt�X������³Z*�
7[=�袏@���>����`��&Mkhd�*!���OG��'z!��/�;:��:g�vr]�d$��`�j\��ѓ��R;ߤn�hHd��qE���z���
�4 I#)�Z'Y��f�t�.��Dn+��Z�>���ɐg�]���U{RH��R� � �b�b�����J�f訅Vq���&�<��} ��.�)l��2�C���|R�|��Il��c����J`!�('�$O�u�Y-�L��[9i���<�C�k��E�[t^���ө?�݆<�aX�@�,G4;�L�m�,�O�$��Q '��>�E�0�ۓ��{���ן\���:�=�b�sM�"��\�^vu�'s�4;�<ZR��wa��D��v��v=�g����҆8��Gb<�fܗ�|`�ï
jJ\��z:���`��QH�*0�:���Ӡ0�h�QY�P��4�?pm�I̅����a,.ͻvWQN]�{���ܰU��S�ꂢ�ui�K�Zr'�|P+ޠH����K�a"���I�_]-И�1n�%@��ع W�	��J���G�����`�
�>�Dj�O�����=_�s�|�̍U�'�Xy|��0�k`qr+	���u ��i��q��e�/C/�B(�`�2ۦϜ��+�۝U��ǡ�Ɖ���"�?ߚ��$�`�x�\>��eL9��j�$mP&G�����Zo���Ƥ
B{4Y��, ��)������yqa4;Y��%ć����ܧ���љ*�!���gJ� ,�ND������q�Ky%��9���"%_/�]	&p��o"�W��lw@�jX�( �g��[��*��u�Y����=Y2T%>�lt}�$.�B��x�}3BW(.�3� ��_�)��sj]���A�ʰĉS��n�0���)��I������p S�2>f��姁�/��A
��$;�q|��D�G�pM|ϴ�N���K���թ 22�1]�m��Ժ�
>0��P�f�A}��1H��y[޽r^*����jb��0�='�s�3Ն��嘭9K�7C����,�2ƿ�h�~H6'��棬VSv�����Eh��;~�ZUݺh�ⴠ�R���KJ�Eu��u�YH�a�%&=���v�M�������[N��R�2�U�����b��;��k��W�Z�V�H��gQ�mW[�LhSc��f���y۫�S�;�ĝ��*'�;���?�wH��jOopVz��y��Tlɷ��N(+s%G~(����?/Lz��_��A03�#}���	��: vzV��.�P(�2�  �S_�2�=1TVl���� 5]O�e|"��q�v�s�tF�N%�:O�����^,�^�0 È�܃���T��=(��C�<�!rq�a�2t�ͪ���C
�)fa� �ޗ��"g=�7�[<����\��t%�xe�Ow��<��xV����M$֛��Z\Ǆ��a���T�A�8B5_C���Q��I���$1~��
tY���S�W İA�.�����i���Z5�I̸��6u4]T� l����0����]�}K�6]�h;G>\�ׅƒ��a�[\�{�g��,苄9��(�͍��4ܢ�`u�� �$�?�9����Oy�hl�\y��u/o>�V�{����>�����'DV�qj���K�Zx��i����{j>}kAх+¹���b=A)�v���q��<>^��(�	R�X��ۈX�6�+f&�1�V{�Rd��/�h�(���\�#̒���pj����t2�VV%Xd�w��Y��:?�ׅ0a�%���7�E*��-�9��ą�Ń�xJ`�z*ӸK$ �����-���u��_��~Q����\������m���?/�%10�Qz�-���3!&�$��ǵ�<+q�Ṯ9���a?P�B���� ��U��,pċ�$�߬i6��x��6ڿ<䚃�J/lvy�C2�X�g�X��|M[����C� ������ ���nǎ{�&��wy�W����]DCv|�5a'�ć"^��j&��
X4�����&��x�R�_��4���%�J�n_@O�9�$�G	e��O`wu@�K�����b�Li&��s��ĳ@P<W#�"��o�����{��a4N�/�c2x�(���ss����ѭ��KO4�B!璩ԡN�s�'kۛe�-*�S��&�׽��l�uf$ET֛L!�_Ln��$)�/��HA`��d�fQ�µ�2�����C&��i�90>��~?��5ގZ9���N�G��V�w����a6T��q��}����<��軓,��*�?���
�U��,`l2y&�	� �g�����r��B��
j}ǭ�k\��/P ��ܮƜĄpR��\H$�]��=�s�$�n�!����Vp�hۓr���o�!���C�X9�q��E�.�h��P�.��x
Xj]R?�<'B���h�ٶ�4��r۰��aq��$�)ɰ/|)0��a�ե���Z]�(����.ΌLhO�s�z��Z_S��v���� %���i��e��-#�A]An:V�g(�%@�[y��^�'�Ւ��N J�Y�eڴ>�1R�!���ԐRq��I��Y��FG!�]Y� �t0	��h��1�Q��q��ʧ��P]'G�%4����ߠS�OA��(`ω�V�|�F�ȕ�򻸇���xޑ���R�F�ڝ2N��ry�>]�l�P��萵�&q/9�H<�i�+��)>�ѓ[ɲ[݊��?�|4��N�Cj܃r�;���q� Q	-���vr��al�P���*���d���i�,S��K���*@;J��o����`L����G��&�<��.^B���µ���Ԥ}3J�J��r�J03ٺ�v��@���d%;��	给���h�˶s�Iצ�j<o`
.ע�5]�ΏJz8\������-�AL�r/�e:�g���cs�â7�C�!X|�-d���n�����}?��[���|,�9����"�� ����_~�/=�������l��Q�~��WW����	;LNX��e׫f�ph�%q��ω�T=*�n҈{��}a��@u�?gd���������#���a{�F��Ϲ$��z��PM3���pREx���B�]e��Ed^}Y�Q2^�ʶ�<;��|���x�c���f�|_T���@8AZ"��<ԑ�X�ꮾ��]1�׻O�O+�c2,̇�p�T\!���N�M��I`!����n0���1�	s]V�� ��]m� f�#X��S"�5� ��h�݇�8U%b "�xק�9a��.����Z~�ϐ`��}�Ui��LGh���e 6�|��J�<!�������a+Zf0'Kˉ#�>a	٣�BM6�5��'ٛ�l��鿮�ͣ��P�?@�W#�J	��]��?q�9L)_ӏZ2E�?�13X^dp����q	I�/Va��0z!>�&���=���g���J�_]w:$��0��K��Bze�� d���=}�tJ��T��b�O@�o?p�L�ن���R)�������i�돆e�H��p���Ģ�'����(�	G�6�/�+�Rč}�֦�7�g]����$��M��i�8��i۲"(�~U��n:�]x'���F�>�,�ñ��i�~A(!<�)F�'�]��͛�|�m��߯06��&�����H6���gv�ZN�M�E�
�ƚ�x��ѱ�z6ae��������m���R���v
��V���������^UW޵����C�{�� 8-Ǫ�1��~�Q�I�>g� N5�������V̝��@��F���g��"�.��|+�`ͭ�pG;k?U���I�SR �F������Wн͠�D�U|���a��Q\��s�׀���v��f����(u"qr�Z0�̣�����L$���x	�Hb�K�Ba<��^�i�F1�����+�<�&2n���c����;_���gV�Ed��WoYo�S�V0�z.�m��oݗ<�^�e�B"�5����g��?ƛ�a���N�^�  �1.d��>�Y��z	��� �_Ȍ�6h"���7T/�B2�JZb���&m��T�v�
�eBL,S��):� ������g��D��<�Z����rh"�c��dq�|�	L!��JƎ���gP��{2"���>�Y�d�u�L���K��q��'�17�s0<������7O��$�f��:l�\]fL��ɧtEa9�I��\mL�m�s`Nu��(i��ً�l���/�����x\��Xd�E��(@0�ԫG������0Әa5�m�.|gNӨjC���pa��=��E͸,�����oޢj�����x,h9����Y�Ht@^0�a6!�{��?���&�a��pbm������6ak���E� �D�&�ɡ�0���̵z�ZS���EdE�#�aɄ��)����Y�V�Re蠕Y�;	���*2����3��������E����~>Ou@���W��&vyҞ�ڀ���8n���Q��Y�,%�G�K�d���`�i�[v�n�&�M�k�M���O���P�8V]���K���/���A� ݈�K]�'ߙ�qeԬ��P=t�q��hL;2�����9@��_o�L�P7	�H�.e��<yS^��*��cGO�:`���L���s&������@c50U���q�s�V��m�V,��q�?ٕu�kcٽs�:}��� o�ƽ���h.$���Ź�O$ӧ���� ��8
(8[�O;�@\qN>(�D爐�-{�D�X�B��! |Aa"O7N����ddX�"��aB�sb��@!v�Lɶ�J)���8n�V4���f�2۷0�IdFk��f��ʅj��hW�~!,RUم�e
֭_���>�Ӿ>�0�-�/z@.Bɲ�-���4ɱ����2�m�����JJ������$�T7փNӺ�YP4"��o
Z�h~<�ʳ�wK#̓��q~�(����ܗ4��+ay�,߶ђ8��<���ۇh���x�/���IU�tS�0����B��4�	o5��YY�-Y���j�KO��`lTY�����h��R��
�lj�#?:��2�9JiZ��J5=R���8���w�A��u�+�DCv@_8��R!-�彐^�>3=fh_q-�c+��
�brvp�9�@���g�1Q�*8M�����	�$6��L)�R��!O�*��Q�
k�j���k�'dUU]�j|B�("�^R�WWI�!��`a��3�"���H貚�G���N�!H�Z)OW��F�s<*q.�Q*{�@J��V3�4X�Á��B��3ۢa�1n1�y����&�cJ,���H��W��eD**w�޸a�{;�S�K@`b�{ws�P��@�����h�	JI�
��V�Æ(O\R��1s��^}ծ4�����V��|eL7���,X �+��[��?KK� ]%����e&�(jL��j6�
F\�p+�Z]~�a��;��FgvC4������$g��C�t��p�����Hpav�T���"ejֳ�Y�i8�Q�􁃱R�VT�	�]�#��.������a����Ʒ�q���+��8R�c-����*x��Ҧ�����\{A6~z�N����bF�Rg]D֚j�����CqX:�!����H5ˢ�g�C=6�o::K8R6�C����e �x2�DW�å�w�YP���	��+��Y��A�e�t;ֈZ�\�2j�=�<�n4� �>
����f�FђY��2)QGrJf?P݉������|Q�&p/���K��4;��>M�2N�[u����^��k�Mv[��XU|b����L[0�%]��½�Ƙ��k^�qN�J\�r�N�����g+��Y4Qn�\ЇAwd�Q�l�#z���h@Q ���t���w��?�Ӕ𙎉v\Ǆ��=��elh�k^4�� ��6\���5ݯd�4��Y����yu�y4���/ *� �!T�L=���	�@���/�U�ȋ��ƋӫI�lj���$d@�,���?�k:��<8��)�X�0�kD������3jJ�J64}ua��:�-�^F
����}��"5f&p��mp&*�`���i� Fb������R����hC�TB��T����T#�S�b}��x�|��m:�ˍn>�����3w�bz9N�b SV�"�r���+Qຨ\����M��Z	R����Үu��]$Iτ�clP�7)sMY)%�.;��x�/B3i�����uܱ]�)A��o�h�Z�vi�J�j�e>���3���0�F�_ U�jŬl���$LQ��ew����֝U�)�<3�a��ض�F{�׬t˖k�����D�6@��� M�|���%�������4��T��"���^^c��R�z7D���Ή�7^�����0��n��=5�c}�_��W{�Q>Tw�TP#>DX��?m��z��[�d����l�uG��j���
]�M��hAٲᱻvwO��ޤ�y�k��[�XK�6��ݯWW90oO��̖�nEv�ruP1	[�� �z�4���ym|D�@d ���UG�m�nC��FK�a �r���у�����1�Z�zSV�t ���+W8��S�}�bpq���&�{k&��L��N}��*��`���Ϗ%��w�U���K3@���"��y�Vm����NWx+���(W��0.���t3��/|�i�Ezo[|p�LD��Q�۠,���<�l����������~I5�͇D�Q�Jly�g��BD�(i+�*=�׈��n�n���F��A��5w�5��^�F��{I ��3�c@71���ɹ��|PN�E�Q�0)���|���5��#�ϨI�?��i�B���H�������r~�?Ղ�n��iE=
%��R��!]��J�]^i�߻XmM1`H Z�A�/:udO㜥�0:��p��<6�.\����[;tT�5�h(X� C}�غ�`���EФ��1]�5��v��Q9a��f�}J���o�X�Kj�����-
���UG�һ�R�j���+ϊ/�p/3A��:��c��bG�������$ic�9eas�Cl�7�����%M|*�(3�v�Fs��$�av��g� "߈�
�)�áF�|$.UP�����H�1�/�d�_ ���������CWR���M�T�1o��Q#x3c��,ۂf����Si�-�`<M��ړl���"���<���a/ۮ���Y�)��xO�.ԍy1�olyHR�dGZ\N���f��3��(��������@�9�z7Ir�6p�)%q��؎TX'�C�{5��k��Ht����~����R�&5��p�:�.�[�)-f��u���u��u�{D�����?Y�!�ۇl�R��me���<��Md�2�n��Xd4�Ȉ���O�^�%p+1�0C�����%a(y�7���o��lV$P��h���:��1��J��	a�L��A��Xu��5�㭊_�["�iY����\>ƽu:�F�R�lQ�yA(�������;]t�a�e��[Ep��ի���>�MY�sQk��{�/X�K�v&�	x���* ����J�ϸ;#��.Ie\����������θj ���	29�s�����c�Fq�{�m�V1��D;A˷o�x���e���T���H]T41���I�d����9�Ǭp�'�xS*��q�'ȯ˙��N�����R� X�)�DW�"G,$�T6y��]�5t���Ժ��H0�9�nB�<3��è�r�?WCֵX��7.�%�ʊ*�ZN;��z���r]1�=�Up����~o��c������]�;�b�S��kJ��֦O�d��5z*��la�5�;_���_d�
��ਨ@��Gj��L���^}�y��\G��Ɍk8�҅�U�8m�RL��������a�����=�x=y�p�;��4p���\����ѷfA��p�x�n�C�@p�<�!����U�j��(Ep8�����V)��Pw$�@8�J*��Ý�yԽ�T]���*���VB���x�Y=M�pZd�LG��U��[4}�H#�`2ֶ�Fa|� z�q�t�>A��,�Z?"Vw��>"
��b/J����{�2�9��	|�3W��J�[2�lT����-_d��R�!�I�R⚌�Χq�|��clV���P��^1d�1�����2n���! ���Hn|� Y:{���f,�ᜠ
b����d�C�I�{�f����mcu��Q����8�+�8�[Q��@V#���D�v���Pя�å�B����q�+}�K��lJ�g�@�����K���\\|���|
U�}a(^�Uͬ���Ը�/.-S�瞇��~�G٫Zz@u�Z=HE������zl��g��lϕ�O��p�ӫ�8�1F�5��=��{W�oH󗩍œי�_7~�z��Df��E�8O9�1`�A�b�h���dt�t�f���M�+�-���uanȄ(�Y����� �Y�s=:1��a(�M�"&9���!�5l�?�ߣ��uh�Ó�榀K�?��Ll���9t]9{�Y�nrn�v�7��NF�^Z�:Kl��u��L�G�gL���n���XxI�����"�[��=LE�yAx��6�y�����Y^č'o��+fA$R�OP+Rmw��6#��!�2�&ݏ�V,_��"s�ב��.���X[�c�f�ʏf&�