��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O��#r#�=�<��/�G��z�nL��u6A[`U1O����K%��g�@�
���I��.�	��q�v\����΃��'rJ����.��J"��ؓ_MG��sG�]��r�5���]�^����$�< �F�u���іQ�^)Jm*�|���j�g�TC��y�h���`g�_�*�ٛ_���j� 7�*����4�t #Z-6 B�x;�ֻH]hE���V]h��Y�\����;�L$�oL��º49R��+�^�1&�q�}��<J	:u���B$5+��@`HO��^a�z�ǎ^Q���⺩�����~�����V�$Oͱk��du˱H��%U�l�q6U`-��MI��>h�P���2�ڡS�2�G��m�)H�w�n_�i����m�����x�3��ecAxa�;��c¶�ZFȤ��AMU�ޕ[��ۦ�m��Ƚ�뇅hs$1��$��Q��;�@6l��xG
��p��t�N4pz�h�2����O�^�����K��g�I�#�(N�̉� X���u(�� t��������qFa�|d�.^;���X�������K+����>��M۔>��H�y��R�8�d|w&�.A��AU6�F�� �c=�|��m�����׬�nL�8�R.Tk8��dϝy�i
4��}�?eP�3�������S���mydTۈ��P�����1g�m�k�VK�ER�H�\��� ��WkpA��P�\"�12�y9Z�V��;@G}˞��X��)/�f!��ΰ]�x��٢��():^� �W�X��t׏�"�[[�Ե��ɖa�eݽILp��Z�(�C�A�ڧ� b4K������4I���:Vn�;o`*Y0��n�!�k;�pj��j,���̅v$�C�2灡iMi!�t��52�Y�2�n�Lǁ�֜�_A>$�rƗ��Ň߯R�2'��d�S!��b`��<E�_s -ͦA��3������ ��f��/��qx�j@xU�kr�Pvnt�9ov�"X�w�����M�S.x5�(���Ot��R�v��tW�����X�D��� O���*���6�qva��UH���ΰjh�	v���z�����9���:Ǹ$H~�j�� ��L����F��\��n�v��#/�%_e3Ed�UG����[H�� (~��[�0|��A	��)��EÌ�]DJ4�X񌖶�J�o�;!���DYոlg
��{M�h8��*�!�Ji�X�:U��4�?�P�8N��,��3ݡ�^�_�X�[���1B�氎��aӜ`P��Y��(E��Kkѷ����`x��PL����{"� ���ȶ���dI�E0XkU�#l/Y�e��O�ܬ,��q!�����,��M,���I�RxZ~�p4O7�����0.���&����}8��v�NtN#�$
�u��=�b{�2E�L{�p��(����5ϻ/D����U���}׺G�V+��虖_b��@Я'��}��I���Uq����W>��ҵf
/�!��)�j��$�P���ndї�w3���&��	�����/�&S��$؇��&��y�W3���cHp�9sx�v�`h�*�� |�6�ݩ�y���<���8�
?$��1}�����P~yl��6cz�b北
����o�<��p���$��mm�R.-��m�6!��e*��mv��
�P������CP��Kc�>���Qg؂��.�9@C�����;��@��+/���၄.�t�ҳ� ��F;=��L�[��5�����~]�]��=G�b�z~��V��"��+�!�4�^���R�LS�w�D����U�KE��(m���O�M�'nS��@Of�p�v��7xd��v4��˟�����ucؿ����;��X�R�l� ���ZF�v 8�R;|w2[�'Mv����O���(?�HO>G�
�Pi���u�����Ν���x� P?r�E�6w���1`�U�m���d8QV9�$�M�3kו�:�Uzլf-{��Ы/w���u�P�<�~A	ѯSҁ��W�)�Ãw��j?-�eʆ�Ѡ��u^��&��3@��q �1?*���j�}@Ŧ���B���A�{1x�4�����ڢ�' ]KV؉\�sE(�}Voѽ�"�>\(���(�l����;^e�B:_'T����	VS'6�(ʞ��7�RҶ��\4��۴�'��Pd�w@���3_�s_58��@�H�� �$6�!��K��Z0��a�+N7al���b.'(;���^t��U`0��v�֊K[�*d�R�����i�f�6��K%�NRg�I�q0���
�~,��ӄ���V[9őò�5pX���\��s�#/�B�UE=eDK����̷cA3�=wV	rp��|�N�%6 I8~l�6x�:?]{<%;<�e����T�3�@PP)13�Y��wS��Ɉ5)�\�Ӱ�+��!�l�:o4��20`Yhƣ|��5�{�"wOQ�gm��T:�JG�[�h���`����5sL�as&��ę&7̍�b�N�ΣԞnm�C�t��ЩD=`bƐۿs<�F��Pz\d���b����N���w����^Vb��Hu�*�m��n4���q���y�l�e�%�:��d�_����w��1C���]�,l�sɜ�.�T;�7/��ς��1��qn�@vP �@e��h@MnY�/��p秬᪹�r&����(Еrf��L�'i�I�^�_�r�OP�+��y�~�;�0�D�߶i�vi!4!,�$b�֜;NW���i-��ď��-�D<Z��a�5J�:��f�$v�d7�v�C�^4��W���14kk�km����,���v�6v���.�����T���'�d�&�Dsx�R�.=��E~.��I~�&ԧ����%�&���ivܐ]�܂�|��9PU:l��?��Y�S�h_�aj�_V�7�%Ͷ�f�o*���H&�|=�n���n�#A���׿_42��D���.S�?�w@,��1�� ��c`2n@M+ӆ�͈�9�OLq�?�̮���l�\��M����\�U�@��*��U�/�ݲڎ�i���U�]�\_�u=�'�+x0�w4a��ט�MH����|r1��Y8|��,dg���Ct�?���~M��q���c��p�HѱN=N5��?kW�p�P'��cp�L�l�� ̫�"����L�K�inS�����D'%|�l���,!�._����2��T�F7\�Kqթ��ߦȊb�E^�K�V����σ���?���(m�͐l��aP�����zy��ȃlÿs1�a�uEɡ������q����MO���&���L�[횠(�^ݾ���'���)u�(����֐q8�)��e �
���ي�%���IF�8 =aW
�� i�ݩ�s8g�Uh��֞ ���H�ț�z_c=肺L SkJ=�}��$T�('�d���o��$���;�0!j��GFL��qf�^��~{V���)���Ja�}�#���=-����X9o�nV� y V�5�vV�Ezn��,����t{��Ϣ&;�5Y���%:^MvO7��H��`{V�
Mm9���CA��oL���Q�zhζT�E�i�h �c�9����y���6!-ܺ�ݬ䫮Q'J�h�.���I�B������ܶd���4�^����Us���
l� �b:���Ђ1��JV��F����2e��I@0tY�N�N��ī`� �0h}���h�3�n�W��̄��T��Ӳ�HK�LH�bX�i*�^VJ����!���a�;�jO���E�mVz�<�v+Ta��׫y����	���)���!r�3��-�ʡ��i���c�
�+����H�JY1ֳ1W�C�x�&���6]����7�����(���+x�?�8p޶=������� Q\�.Ϛz[>�<x�>�D�s�і���M9�y����4�2PH������D(7OQ��^ld>�+����޵n�W�8Guw ��) <Եz�wBԆ���Q p��߫����}���V��Uf����k�� �)�b�uȪn�R� �����I�,��vs�F���̈́S5��,~�K��q/����H�����-x��qV��>�%�(<�v�Cq�yNPކ�f���G6ův��+60�]=mMg;ꧾu��X�ђ�*N�#�c���Z�7�m#rtY����(	v�&�:&��{����Yބ�OOf���^�XҌ�/����*�xܦ-����!��ӕ*>|�<
J�����CI���va�v5��
�0ۇ\��w�4* �)��yG$㜕X��kc����
�=��N����	��4W��z����ƾR�J��^��2;���Z�W2%d�Y��?{`�T���,�r�ۊ�ukh��͢k� `��Tm���͢g�����PK�H�K�:��2��($j�+��<�40�I��n)�`MAB=o���N�6p�hR=.���2�U�:�j�v��ꆾK�%�7ȶ��'�!1������lNb/4����.3��;��5Sy��O��9����X�}%h�ǂ�?J�Pe��D��H������g��'3;y&���[����ב?��� ���H�e��#��l��q�����݇�x��+�cM�n��EB���E] ����*lX�Q+ [���p{�:C�
�ը��=�\��婭";���7f�/_��"��Z�Lh>�	�% ����IR[���M t*xZE���"���z[�����ţ�~  ����3.ƉĜ��xU.s��nYa�;���i����c/G�F�BL�h]�?��-���k��%�K�=�mH��,�Q� b��?A8��y}������ԅ�P6��R�E�xS����>����$Ϛ�S�Ö@H�ͥ���r� ���D��1�����%,��_}�E�ā��(<N@~T�f�E�<{�26���
�$�wMO��QeÐ.�Z+̿��d.�+�_̚/T'��<h��G��d�^DJ���M�m��	�Ͼ��<���x5oo��=&{�h�(�H�CnPZ�Ē�@Ndې=��	陸�'�; ��$����[߻��������n����7�@N�Z�ML�B@PO�	�zI����Q�b���=ؼ�㛠�?�QJ��;H�+Do9��D���1��2,��Ѓb�nB@��T5'��I���H����y����!{�0*��Qɒ.�}�-�����@�	�������떳s�ϖ����v<�,�GYh�g!tq�pτ�^�73˽�
��L�Vh��ʘX%�H� �a
u�'(u������aE	�Ω�Ppsr�b��L]$/6!�z_�7������A�$/
����Z����\�������:e2��Oҏeݴ�ф7�a���saJ>��C�<)�֎�cǻ���@�����p{��=�Xg�C_�]��b����- �̜�0!��Nn�䫯��(>�]������L�}��Ɗ�2��a�c�[�� !O,iwل�e{ �t�W?�H�y�<���W�L�!�Gn5F�T���b�3.�b�7�bq;\�7�7Tp1o��5�|��;V�7g.)p3�k�0)�
��+���4��t%�$|�A(0n��s�T�@�/�ϡ�W%���-������J�UCس:m�����0���4 ���I�����^�~�o�Y�XK}��+��Ǉ���_�0�LI���rF��V�9����K�\�'7d\�KfsJ�yw9~:��}�̕ijc��[ژ��:�Y�]6����@�o��L>�pho-P����W�u�MiD�>�ρ�P�B�}V�A��+aW���no�\H��鹺-!��(U��^5r_�nʜ����|'����o�����]ȳ2�KlQ۽��7��?��~7�[Y��[_k���U�Y�J�VW�)�"�����d�w���*rQ�X�IDrm�u4w����E�+RGUQ�m�C�B�4h��k;�/��J'�X7�W�����}���<����Bz��;���l	������_��`>�۰�Z���䣈` ��%�%�E\�|�V^+�t�%�p��V�"��;�0V���H?9������,�@KY���^�&�G��$��G��<X��r- i���qq���K�u^���MAPD���6H���7k��Y~��4D�0\�n�0�Մ���q/oG2���_fa,x0mrvў�&����{!u����7o`|��G�M��pь�6�m���<7N>��}�YR�W�iJ>�
�R���.c�s(� ��X�Aa��[Qc +�Z:_��^�8��X!e�/kk�(X�RաHX���ˍXn� �f��'�,�����їC�����K�.T���T���}��iM��#�����O(`��<�oY ���y���u�J�o������t�
��t\�v�+�uE�f!9�$�L���Vl�I7�FA�..۫XA��0��F�2��F�c���.�D-@��z�=Ep�����MG. ���a�t�\�
���>��g��X� @5sh��_��n��K(����^�S�{�h�O�MN�ʱ? ��'r�r�_��
�)4 �۪��m�r����τ{��Y�0+��muno���A�a{��޺�=���y5�?�v�P���(�-Q�2(��9�J�d�nǺׄ{?$}sx�e����뢎wSq��o��J�W&+ۿ�ƣ�m�-�����aBȨ
:�нӤ�fu��J�vz��/�h����WR�%x���h�h�q�G��;MV�K�VM>�h]�B�\x�Y��хL�f������~�Wi��=i�\w���ހ���j���'=��U+5���+����[̄f�Y�l���x%